`define FORCE_NO_INSTANTIATE_TM1638_BOARD_CONTROLLER_MODULE
`include "../tang_nano_4k_hdmi_tm1638/board_specific_top.sv"
