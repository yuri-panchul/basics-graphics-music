`include "../nexys_a7_100/board_specific_top.sv"
