`define USE_LCD_800_480
`include "../tang_nano_20k_lcd_480_272_tm1638/board_specific_top.sv"
