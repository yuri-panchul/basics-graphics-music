`include "config.svh"

module tb;

    testbench i_tb ();

endmodule
