`define ALINX_AX4010
`include "../saylinx/board_specific_top.sv"
