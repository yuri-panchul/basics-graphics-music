`define FORCE_NO_INSTANTIATE_TM1638_BOARD_CONTROLLER_MODULE
`define USE_LCD_480_272_ML6485
`include "../tang_nano_9k_lcd_480_272_tm1638/board_specific_top.sv"
