`define USE_HACKATHON_TOP
`include "../tang_nano_9k_lcd_480_272_tm1638/board_specific_top.sv"
