`define VGA666_BOARD
`include "../de0_nano_vga_pmod/board_specific_top.sv"
