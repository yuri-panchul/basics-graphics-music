`define USE_DIGILENT_PMOD_MIC3
`include "../omdazz/board_specific_top.sv"
