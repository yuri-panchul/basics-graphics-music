// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=261.63Hz, Fs=48828Hz, 16-bit, Volume 100%

module table_48828_C
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 47;

    always_comb
        case (x)
         0: y = 16'b0000000000000000;
         1: y = 16'b0000001111011001;
         2: y = 16'b0000011110110010;
         3: y = 16'b0000101110001000;
         4: y = 16'b0000111101011011;
         5: y = 16'b0001001100101001;
         6: y = 16'b0001011011110010;
         7: y = 16'b0001101010110101;
         8: y = 16'b0001111001110000;
         9: y = 16'b0010001000100010;
        10: y = 16'b0010010111001010;
        11: y = 16'b0010100101101000;
        12: y = 16'b0010110011111001;
        13: y = 16'b0011000001111110;
        14: y = 16'b0011001111110101;
        15: y = 16'b0011011101011101;
        16: y = 16'b0011101010110110;
        17: y = 16'b0011110111111101;
        18: y = 16'b0100000100110011;
        19: y = 16'b0100010001010110;
        20: y = 16'b0100011101100110;
        21: y = 16'b0100101001100001;
        22: y = 16'b0100110101000111;
        23: y = 16'b0101000000010111;
        24: y = 16'b0101001011010000;
        25: y = 16'b0101010101110001;
        26: y = 16'b0101011111111010;
        27: y = 16'b0101101001101001;
        28: y = 16'b0101110010111111;
        29: y = 16'b0101111011111010;
        30: y = 16'b0110000100011011;
        31: y = 16'b0110001100011111;
        32: y = 16'b0110010100000111;
        33: y = 16'b0110011011010010;
        34: y = 16'b0110100010000000;
        35: y = 16'b0110101000010000;
        36: y = 16'b0110101110000001;
        37: y = 16'b0110110011010100;
        38: y = 16'b0110111000001000;
        39: y = 16'b0110111100011100;
        40: y = 16'b0111000000010001;
        41: y = 16'b0111000011100101;
        42: y = 16'b0111000110011001;
        43: y = 16'b0111001000101101;
        44: y = 16'b0111001010100000;
        45: y = 16'b0111001011110010;
        46: y = 16'b0111001100100100;
        47: y = 16'b0111001100110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=277.18Hz, Fs=48828Hz, 16-bit, Volume 100%

module table_48828_Cs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 44;

    always_comb
        case (x)
         0: y = 16'b0000000000000000;
         1: y = 16'b0000010000011101;
         2: y = 16'b0000100000111000;
         3: y = 16'b0000110001010001;
         4: y = 16'b0001000001100101;
         5: y = 16'b0001010001110100;
         6: y = 16'b0001100001111101;
         7: y = 16'b0001110001111110;
         8: y = 16'b0010000001110101;
         9: y = 16'b0010010001100010;
        10: y = 16'b0010100001000010;
        11: y = 16'b0010110000010110;
        12: y = 16'b0010111111011011;
        13: y = 16'b0011001110010001;
        14: y = 16'b0011011100110110;
        15: y = 16'b0011101011001001;
        16: y = 16'b0011111001001001;
        17: y = 16'b0100000110110100;
        18: y = 16'b0100010100001010;
        19: y = 16'b0100100001001001;
        20: y = 16'b0100101101110001;
        21: y = 16'b0100111010000000;
        22: y = 16'b0101000101110110;
        23: y = 16'b0101010001010001;
        24: y = 16'b0101011100010001;
        25: y = 16'b0101100110110100;
        26: y = 16'b0101110000111010;
        27: y = 16'b0101111010100001;
        28: y = 16'b0110000011101010;
        29: y = 16'b0110001100010100;
        30: y = 16'b0110010100011101;
        31: y = 16'b0110011100000100;
        32: y = 16'b0110100011001011;
        33: y = 16'b0110101001101111;
        34: y = 16'b0110101111110001;
        35: y = 16'b0110110101001111;
        36: y = 16'b0110111010001001;
        37: y = 16'b0110111110100000;
        38: y = 16'b0111000010010010;
        39: y = 16'b0111000101011111;
        40: y = 16'b0111001000001000;
        41: y = 16'b0111001010001011;
        42: y = 16'b0111001011101001;
        43: y = 16'b0111001100100001;
        44: y = 16'b0111001100110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=293.66Hz, Fs=48828Hz, 16-bit, Volume 100%

module table_48828_D
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 42;

    always_comb
        case (x)
         0: y = 16'b0000000000000000;
         1: y = 16'b0000010001001111;
         2: y = 16'b0000100010011100;
         3: y = 16'b0000110011100110;
         4: y = 16'b0001000100101100;
         5: y = 16'b0001010101101011;
         6: y = 16'b0001100110100011;
         7: y = 16'b0001110111010001;
         8: y = 16'b0010000111110101;
         9: y = 16'b0010011000001101;
        10: y = 16'b0010101000010111;
        11: y = 16'b0010111000010010;
        12: y = 16'b0011000111111100;
        13: y = 16'b0011010111010101;
        14: y = 16'b0011100110011010;
        15: y = 16'b0011110101001011;
        16: y = 16'b0100000011100101;
        17: y = 16'b0100010001101001;
        18: y = 16'b0100011111010100;
        19: y = 16'b0100101100100101;
        20: y = 16'b0100111001011100;
        21: y = 16'b0101000101110110;
        22: y = 16'b0101010001110011;
        23: y = 16'b0101011101010010;
        24: y = 16'b0101101000010010;
        25: y = 16'b0101110010110001;
        26: y = 16'b0101111100101111;
        27: y = 16'b0110000110001100;
        28: y = 16'b0110001111000101;
        29: y = 16'b0110010111011010;
        30: y = 16'b0110011111001011;
        31: y = 16'b0110100110010111;
        32: y = 16'b0110101100111101;
        33: y = 16'b0110110010111101;
        34: y = 16'b0110111000010110;
        35: y = 16'b0110111101000111;
        36: y = 16'b0111000001010001;
        37: y = 16'b0111000100110010;
        38: y = 16'b0111000111101011;
        39: y = 16'b0111001001111011;
        40: y = 16'b0111001011100010;
        41: y = 16'b0111001100011111;
        42: y = 16'b0111001100110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=311.13Hz, Fs=48828Hz, 16-bit, Volume 100%

module table_48828_Ds
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 39;

    always_comb
        case (x)
         0: y = 16'b0000000000000000;
         1: y = 16'b0000010010100100;
         2: y = 16'b0000100101000101;
         3: y = 16'b0000110111100011;
         4: y = 16'b0001001001111011;
         5: y = 16'b0001011100001011;
         6: y = 16'b0001101110010010;
         7: y = 16'b0010000000001101;
         8: y = 16'b0010010001111011;
         9: y = 16'b0010100011011010;
        10: y = 16'b0010110100101000;
        11: y = 16'b0011000101100011;
        12: y = 16'b0011010110001010;
        13: y = 16'b0011100110011010;
        14: y = 16'b0011110110010010;
        15: y = 16'b0100000101110001;
        16: y = 16'b0100010100110101;
        17: y = 16'b0100100011011100;
        18: y = 16'b0100110001100101;
        19: y = 16'b0100111111001110;
        20: y = 16'b0101001100010110;
        21: y = 16'b0101011000111011;
        22: y = 16'b0101100100111101;
        23: y = 16'b0101110000011001;
        24: y = 16'b0101111011001111;
        25: y = 16'b0110000101011110;
        26: y = 16'b0110001111000101;
        27: y = 16'b0110011000000010;
        28: y = 16'b0110100000010101;
        29: y = 16'b0110100111111100;
        30: y = 16'b0110101110110111;
        31: y = 16'b0110110101000110;
        32: y = 16'b0110111010101000;
        33: y = 16'b0110111111011011;
        34: y = 16'b0111000011100000;
        35: y = 16'b0111000110110110;
        36: y = 16'b0111001001011101;
        37: y = 16'b0111001011010100;
        38: y = 16'b0111001100011100;
        39: y = 16'b0111001100110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=329.63Hz, Fs=48828Hz, 16-bit, Volume 100%

module table_48828_E
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 37;

    always_comb
        case (x)
         0: y = 16'b0000000000000000;
         1: y = 16'b0000010011100100;
         2: y = 16'b0000100111000101;
         3: y = 16'b0000111010100010;
         4: y = 16'b0001001101111000;
         5: y = 16'b0001100001000101;
         6: y = 16'b0001110100000111;
         7: y = 16'b0010000110111100;
         8: y = 16'b0010011001100001;
         9: y = 16'b0010101011110100;
        10: y = 16'b0010111101110100;
        11: y = 16'b0011001111011101;
        12: y = 16'b0011100000101111;
        13: y = 16'b0011110001100111;
        14: y = 16'b0100000010000011;
        15: y = 16'b0100010010000001;
        16: y = 16'b0100100001011111;
        17: y = 16'b0100110000011101;
        18: y = 16'b0100111110110111;
        19: y = 16'b0101001100101100;
        20: y = 16'b0101011001111011;
        21: y = 16'b0101100110100010;
        22: y = 16'b0101110010011111;
        23: y = 16'b0101111101110010;
        24: y = 16'b0110001000011001;
        25: y = 16'b0110010010010011;
        26: y = 16'b0110011011011110;
        27: y = 16'b0110100011111010;
        28: y = 16'b0110101011100101;
        29: y = 16'b0110110010011111;
        30: y = 16'b0110111000100111;
        31: y = 16'b0110111101111100;
        32: y = 16'b0111000010011110;
        33: y = 16'b0111000110001100;
        34: y = 16'b0111001001000101;
        35: y = 16'b0111001011001010;
        36: y = 16'b0111001100011001;
        37: y = 16'b0111001100110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=349.23Hz, Fs=48828Hz, 16-bit, Volume 100%

module table_48828_F
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 35;

    always_comb
        case (x)
         0: y = 16'b0000000000000000;
         1: y = 16'b0000010100101011;
         2: y = 16'b0000101001010100;
         3: y = 16'b0000111101110111;
         4: y = 16'b0001010010010010;
         5: y = 16'b0001100110100011;
         6: y = 16'b0001111010100110;
         7: y = 16'b0010001110011010;
         8: y = 16'b0010100001111011;
         9: y = 16'b0010110101000111;
        10: y = 16'b0011000111111100;
        11: y = 16'b0011011010010111;
        12: y = 16'b0011101100010110;
        13: y = 16'b0011111101110111;
        14: y = 16'b0100001110110111;
        15: y = 16'b0100011111010100;
        16: y = 16'b0100101111001100;
        17: y = 16'b0100111110011101;
        18: y = 16'b0101001101000101;
        19: y = 16'b0101011011000010;
        20: y = 16'b0101101000010010;
        21: y = 16'b0101110100110100;
        22: y = 16'b0110000000100101;
        23: y = 16'b0110001011100101;
        24: y = 16'b0110010101110011;
        25: y = 16'b0110011111001011;
        26: y = 16'b0110100111101111;
        27: y = 16'b0110101111011011;
        28: y = 16'b0110110110010001;
        29: y = 16'b0110111100001101;
        30: y = 16'b0111000001010001;
        31: y = 16'b0111000101011010;
        32: y = 16'b0111001000101001;
        33: y = 16'b0111001010111101;
        34: y = 16'b0111001100010110;
        35: y = 16'b0111001100110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=369.99Hz, Fs=48828Hz, 16-bit, Volume 100%

module table_48828_Fs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 33;

    always_comb
        case (x)
         0: y = 16'b0000000000000000;
         1: y = 16'b0000010101111011;
         2: y = 16'b0000101011110011;
         3: y = 16'b0001000001100101;
         4: y = 16'b0001010111001101;
         5: y = 16'b0001101100101001;
         6: y = 16'b0010000001110101;
         7: y = 16'b0010010110101110;
         8: y = 16'b0010101011010001;
         9: y = 16'b0010111111011011;
        10: y = 16'b0011010011001010;
        11: y = 16'b0011100110011010;
        12: y = 16'b0011111001001001;
        13: y = 16'b0100001011010011;
        14: y = 16'b0100011100110111;
        15: y = 16'b0100101101110001;
        16: y = 16'b0100111110000000;
        17: y = 16'b0101001101100000;
        18: y = 16'b0101011100010001;
        19: y = 16'b0101101010001110;
        20: y = 16'b0101110111010111;
        21: y = 16'b0110000011101010;
        22: y = 16'b0110001111000101;
        23: y = 16'b0110011001100110;
        24: y = 16'b0110100011001011;
        25: y = 16'b0110101011110011;
        26: y = 16'b0110110011011110;
        27: y = 16'b0110111010001001;
        28: y = 16'b0110111111110101;
        29: y = 16'b0111000100011111;
        30: y = 16'b0111001000001000;
        31: y = 16'b0111001010101110;
        32: y = 16'b0111001100010011;
        33: y = 16'b0111001100110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=392.0Hz, Fs=48828Hz, 16-bit, Volume 100%

module table_48828_G
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 31;

    always_comb
        case (x)
         0: y = 16'b0000000000000000;
         1: y = 16'b0000010111010110;
         2: y = 16'b0000101110101000;
         3: y = 16'b0001000101110010;
         4: y = 16'b0001011100110001;
         5: y = 16'b0001110011100000;
         6: y = 16'b0010001001111101;
         7: y = 16'b0010100000000011;
         8: y = 16'b0010110101101110;
         9: y = 16'b0011001010111100;
        10: y = 16'b0011011111101001;
        11: y = 16'b0011110011110000;
        12: y = 16'b0100000111010000;
        13: y = 16'b0100011010000100;
        14: y = 16'b0100101100001010;
        15: y = 16'b0100111101011111;
        16: y = 16'b0101001110000000;
        17: y = 16'b0101011101101001;
        18: y = 16'b0101101100011010;
        19: y = 16'b0101111010001110;
        20: y = 16'b0110000111000100;
        21: y = 16'b0110010010111010;
        22: y = 16'b0110011101101110;
        23: y = 16'b0110100111011110;
        24: y = 16'b0110110000001000;
        25: y = 16'b0110110111101011;
        26: y = 16'b0110111110000111;
        27: y = 16'b0111000011011000;
        28: y = 16'b0111000111100000;
        29: y = 16'b0111001010011101;
        30: y = 16'b0111001100001110;
        31: y = 16'b0111001100110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=415.3Hz, Fs=48828Hz, 16-bit, Volume 100%

module table_48828_Gs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 29;

    always_comb
        case (x)
         0: y = 16'b0000000000000000;
         1: y = 16'b0000011000111101;
         2: y = 16'b0000110001110101;
         3: y = 16'b0001001010100011;
         4: y = 16'b0001100011000100;
         5: y = 16'b0001111011010010;
         6: y = 16'b0010010011001001;
         7: y = 16'b0010101010100100;
         8: y = 16'b0011000001011111;
         9: y = 16'b0011010111110110;
        10: y = 16'b0011101101100101;
        11: y = 16'b0100000010100111;
        12: y = 16'b0100010110111000;
        13: y = 16'b0100101010010101;
        14: y = 16'b0100111100111010;
        15: y = 16'b0101001110100011;
        16: y = 16'b0101011111001110;
        17: y = 16'b0101101110110110;
        18: y = 16'b0101111101011010;
        19: y = 16'b0110001010110110;
        20: y = 16'b0110010111001001;
        21: y = 16'b0110100010001110;
        22: y = 16'b0110101100000101;
        23: y = 16'b0110110100101100;
        24: y = 16'b0110111100000001;
        25: y = 16'b0111000010000010;
        26: y = 16'b0111000110101111;
        27: y = 16'b0111001010000111;
        28: y = 16'b0111001100001001;
        29: y = 16'b0111001100110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=440.0Hz, Fs=48828Hz, 16-bit, Volume 100%

module table_48828_A
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 28;

    always_comb
        case (x)
         0: y = 16'b0000000000000000;
         1: y = 16'b0000011001110110;
         2: y = 16'b0000110011100110;
         3: y = 16'b0001001101001100;
         4: y = 16'b0001100110100011;
         5: y = 16'b0001111111100100;
         6: y = 16'b0010011000001101;
         7: y = 16'b0010110000010110;
         8: y = 16'b0011000111111100;
         9: y = 16'b0011011110111010;
        10: y = 16'b0011110101001011;
        11: y = 16'b0100001010101010;
        12: y = 16'b0100011111010100;
        13: y = 16'b0100110011000100;
        14: y = 16'b0101000101110110;
        15: y = 16'b0101010111100110;
        16: y = 16'b0101101000010010;
        17: y = 16'b0101110111110101;
        18: y = 16'b0110000110001100;
        19: y = 16'b0110010011010100;
        20: y = 16'b0110011111001011;
        21: y = 16'b0110101001101111;
        22: y = 16'b0110110010111101;
        23: y = 16'b0110111010110011;
        24: y = 16'b0111000001010001;
        25: y = 16'b0111000110010011;
        26: y = 16'b0111001001111011;
        27: y = 16'b0111001100000110;
        28: y = 16'b0111001100110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=466.16Hz, Fs=48828Hz, 16-bit, Volume 100%

module table_48828_As
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 26;

    always_comb
        case (x)
         0: y = 16'b0000000000000000;
         1: y = 16'b0000011011110101;
         2: y = 16'b0000110111100011;
         3: y = 16'b0001010011000100;
         4: y = 16'b0001101110010010;
         5: y = 16'b0010001001000110;
         6: y = 16'b0010100011011010;
         7: y = 16'b0010111101001000;
         8: y = 16'b0011010110001010;
         9: y = 16'b0011101110011001;
        10: y = 16'b0100000101110001;
        11: y = 16'b0100011100001100;
        12: y = 16'b0100110001100101;
        13: y = 16'b0101000101110110;
        14: y = 16'b0101011000111011;
        15: y = 16'b0101101010110000;
        16: y = 16'b0101111011001111;
        17: y = 16'b0110001010010111;
        18: y = 16'b0110011000000010;
        19: y = 16'b0110100100001110;
        20: y = 16'b0110101110110111;
        21: y = 16'b0110110111111101;
        22: y = 16'b0110111111011011;
        23: y = 16'b0111000101010001;
        24: y = 16'b0111001001011101;
        25: y = 16'b0111001011111110;
        26: y = 16'b0111001100110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=493.88Hz, Fs=48828Hz, 16-bit, Volume 100%

module table_48828_B
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 25;

    always_comb
        case (x)
         0: y = 16'b0000000000000000;
         1: y = 16'b0000011100111100;
         2: y = 16'b0000111001110000;
         3: y = 16'b0001010110010110;
         4: y = 16'b0001110010100110;
         5: y = 16'b0010001110011010;
         6: y = 16'b0010101001101001;
         7: y = 16'b0011000100001101;
         8: y = 16'b0011011110000000;
         9: y = 16'b0011110110111011;
        10: y = 16'b0100001110110111;
        11: y = 16'b0100100101101111;
        12: y = 16'b0100111011011101;
        13: y = 16'b0101001111111011;
        14: y = 16'b0101100011000100;
        15: y = 16'b0101110100110100;
        16: y = 16'b0110000101000101;
        17: y = 16'b0110010011110100;
        18: y = 16'b0110100000111101;
        19: y = 16'b0110101100011101;
        20: y = 16'b0110110110010001;
        21: y = 16'b0110111110010101;
        22: y = 16'b0111000100101010;
        23: y = 16'b0111001001001011;
        24: y = 16'b0111001011111010;
        25: y = 16'b0111001100110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=261.63Hz, Fs=64453Hz, 16-bit, Volume 100%

module table_64453_C
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 62;

    always_comb
        case (x)
         0: y = 16'b0000000000000000;
         1: y = 16'b0000001011101011;
         2: y = 16'b0000010111010110;
         3: y = 16'b0000100010111111;
         4: y = 16'b0000101110101000;
         5: y = 16'b0000111010001110;
         6: y = 16'b0001000101110010;
         7: y = 16'b0001010001010011;
         8: y = 16'b0001011100110001;
         9: y = 16'b0001101000001011;
        10: y = 16'b0001110011100000;
        11: y = 16'b0001111110110001;
        12: y = 16'b0010001001111101;
        13: y = 16'b0010010101000011;
        14: y = 16'b0010100000000011;
        15: y = 16'b0010101010111100;
        16: y = 16'b0010110101101110;
        17: y = 16'b0011000000011001;
        18: y = 16'b0011001010111100;
        19: y = 16'b0011010101010111;
        20: y = 16'b0011011111101001;
        21: y = 16'b0011101001110001;
        22: y = 16'b0011110011110000;
        23: y = 16'b0011111101100101;
        24: y = 16'b0100000111010000;
        25: y = 16'b0100010000110000;
        26: y = 16'b0100011010000100;
        27: y = 16'b0100100011001101;
        28: y = 16'b0100101100001010;
        29: y = 16'b0100110100111011;
        30: y = 16'b0100111101011111;
        31: y = 16'b0101000101110110;
        32: y = 16'b0101001110000000;
        33: y = 16'b0101010101111011;
        34: y = 16'b0101011101101001;
        35: y = 16'b0101100101001001;
        36: y = 16'b0101101100011010;
        37: y = 16'b0101110011011011;
        38: y = 16'b0101111010001110;
        39: y = 16'b0110000000110001;
        40: y = 16'b0110000111000100;
        41: y = 16'b0110001101000111;
        42: y = 16'b0110010010111010;
        43: y = 16'b0110011000011101;
        44: y = 16'b0110011101101110;
        45: y = 16'b0110100010101111;
        46: y = 16'b0110100111011110;
        47: y = 16'b0110101011111100;
        48: y = 16'b0110110000001000;
        49: y = 16'b0110110100000011;
        50: y = 16'b0110110111101011;
        51: y = 16'b0110111011000010;
        52: y = 16'b0110111110000111;
        53: y = 16'b0111000000111001;
        54: y = 16'b0111000011011000;
        55: y = 16'b0111000101100101;
        56: y = 16'b0111000111100000;
        57: y = 16'b0111001001001000;
        58: y = 16'b0111001010011101;
        59: y = 16'b0111001011011111;
        60: y = 16'b0111001100001110;
        61: y = 16'b0111001100101011;
        62: y = 16'b0111001100110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=277.18Hz, Fs=64453Hz, 16-bit, Volume 100%

module table_64453_Cs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 58;

    always_comb
        case (x)
         0: y = 16'b0000000000000000;
         1: y = 16'b0000001100011111;
         2: y = 16'b0000011000111101;
         3: y = 16'b0000100101011010;
         4: y = 16'b0000110001110101;
         5: y = 16'b0000111110001101;
         6: y = 16'b0001001010100011;
         7: y = 16'b0001010110110110;
         8: y = 16'b0001100011000100;
         9: y = 16'b0001101111001110;
        10: y = 16'b0001111011010010;
        11: y = 16'b0010000111010001;
        12: y = 16'b0010010011001001;
        13: y = 16'b0010011110111010;
        14: y = 16'b0010101010100100;
        15: y = 16'b0010110110000110;
        16: y = 16'b0011000001011111;
        17: y = 16'b0011001100110000;
        18: y = 16'b0011010111110110;
        19: y = 16'b0011100010110011;
        20: y = 16'b0011101101100101;
        21: y = 16'b0011111000001011;
        22: y = 16'b0100000010100111;
        23: y = 16'b0100001100110101;
        24: y = 16'b0100010110111000;
        25: y = 16'b0100100000101101;
        26: y = 16'b0100101010010101;
        27: y = 16'b0100110011101110;
        28: y = 16'b0100111100111010;
        29: y = 16'b0101000101110110;
        30: y = 16'b0101001110100011;
        31: y = 16'b0101010111000000;
        32: y = 16'b0101011111001110;
        33: y = 16'b0101100111001010;
        34: y = 16'b0101101110110110;
        35: y = 16'b0101110110010001;
        36: y = 16'b0101111101011010;
        37: y = 16'b0110000100010001;
        38: y = 16'b0110001010110110;
        39: y = 16'b0110010001001001;
        40: y = 16'b0110010111001001;
        41: y = 16'b0110011100110101;
        42: y = 16'b0110100010001110;
        43: y = 16'b0110100111010100;
        44: y = 16'b0110101100000101;
        45: y = 16'b0110110000100011;
        46: y = 16'b0110110100101100;
        47: y = 16'b0110111000100001;
        48: y = 16'b0110111100000001;
        49: y = 16'b0110111111001100;
        50: y = 16'b0111000010000010;
        51: y = 16'b0111000100100100;
        52: y = 16'b0111000110101111;
        53: y = 16'b0111001000100110;
        54: y = 16'b0111001010000111;
        55: y = 16'b0111001011010011;
        56: y = 16'b0111001100001001;
        57: y = 16'b0111001100101001;
        58: y = 16'b0111001100110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=293.66Hz, Fs=64453Hz, 16-bit, Volume 100%

module table_64453_D
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 55;

    always_comb
        case (x)
         0: y = 16'b0000000000000000;
         1: y = 16'b0000001101001010;
         2: y = 16'b0000011010010100;
         3: y = 16'b0000100111011100;
         4: y = 16'b0000110100100010;
         5: y = 16'b0001000001100101;
         6: y = 16'b0001001110100101;
         7: y = 16'b0001011011100001;
         8: y = 16'b0001101000011000;
         9: y = 16'b0001110101001001;
        10: y = 16'b0010000001110101;
        11: y = 16'b0010001110011010;
        12: y = 16'b0010011010110111;
        13: y = 16'b0010100111001100;
        14: y = 16'b0010110011011000;
        15: y = 16'b0010111111011011;
        16: y = 16'b0011001011010100;
        17: y = 16'b0011010111000011;
        18: y = 16'b0011100010100110;
        19: y = 16'b0011101101111110;
        20: y = 16'b0011111001001001;
        21: y = 16'b0100000100000111;
        22: y = 16'b0100001110110111;
        23: y = 16'b0100011001011001;
        24: y = 16'b0100100011101101;
        25: y = 16'b0100101101110001;
        26: y = 16'b0100110111100110;
        27: y = 16'b0101000001001010;
        28: y = 16'b0101001010011110;
        29: y = 16'b0101010011100000;
        30: y = 16'b0101011100010001;
        31: y = 16'b0101100100101111;
        32: y = 16'b0101101100111011;
        33: y = 16'b0101110100110100;
        34: y = 16'b0101111100011001;
        35: y = 16'b0110000011101010;
        36: y = 16'b0110001010100111;
        37: y = 16'b0110010001010000;
        38: y = 16'b0110010111100100;
        39: y = 16'b0110011101100010;
        40: y = 16'b0110100011001011;
        41: y = 16'b0110101000011110;
        42: y = 16'b0110101101011011;
        43: y = 16'b0110110010000001;
        44: y = 16'b0110110110010001;
        45: y = 16'b0110111010001001;
        46: y = 16'b0110111101101011;
        47: y = 16'b0111000000110110;
        48: y = 16'b0111000011101001;
        49: y = 16'b0111000110000100;
        50: y = 16'b0111001000001000;
        51: y = 16'b0111001001110100;
        52: y = 16'b0111001011001000;
        53: y = 16'b0111001100000100;
        54: y = 16'b0111001100101000;
        55: y = 16'b0111001100110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=311.13Hz, Fs=64453Hz, 16-bit, Volume 100%

module table_64453_Ds
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 52;

    always_comb
        case (x)
         0: y = 16'b0000000000000000;
         1: y = 16'b0000001101111011;
         2: y = 16'b0000011011110101;
         3: y = 16'b0000101001101101;
         4: y = 16'b0000110111100011;
         5: y = 16'b0001000101010101;
         6: y = 16'b0001010011000100;
         7: y = 16'b0001100000101110;
         8: y = 16'b0001101110010010;
         9: y = 16'b0001111011110000;
        10: y = 16'b0010001001000110;
        11: y = 16'b0010010110010100;
        12: y = 16'b0010100011011010;
        13: y = 16'b0010110000010110;
        14: y = 16'b0010111101001000;
        15: y = 16'b0011001001101111;
        16: y = 16'b0011010110001010;
        17: y = 16'b0011100010011000;
        18: y = 16'b0011101110011001;
        19: y = 16'b0011111010001101;
        20: y = 16'b0100000101110001;
        21: y = 16'b0100010001000111;
        22: y = 16'b0100011100001100;
        23: y = 16'b0100100111000001;
        24: y = 16'b0100110001100101;
        25: y = 16'b0100111011110111;
        26: y = 16'b0101000101110110;
        27: y = 16'b0101001111100010;
        28: y = 16'b0101011000111011;
        29: y = 16'b0101100010000000;
        30: y = 16'b0101101010110000;
        31: y = 16'b0101110011001010;
        32: y = 16'b0101111011001111;
        33: y = 16'b0110000010111110;
        34: y = 16'b0110001010010111;
        35: y = 16'b0110010001011000;
        36: y = 16'b0110011000000010;
        37: y = 16'b0110011110010100;
        38: y = 16'b0110100100001110;
        39: y = 16'b0110101001101111;
        40: y = 16'b0110101110110111;
        41: y = 16'b0110110011100111;
        42: y = 16'b0110110111111101;
        43: y = 16'b0110111011111001;
        44: y = 16'b0110111111011011;
        45: y = 16'b0111000010100011;
        46: y = 16'b0111000101010001;
        47: y = 16'b0111000111100100;
        48: y = 16'b0111001001011101;
        49: y = 16'b0111001010111011;
        50: y = 16'b0111001011111110;
        51: y = 16'b0111001100100111;
        52: y = 16'b0111001100110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=329.63Hz, Fs=64453Hz, 16-bit, Volume 100%

module table_64453_E
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 49;

    always_comb
        case (x)
         0: y = 16'b0000000000000000;
         1: y = 16'b0000001110110001;
         2: y = 16'b0000011101100010;
         3: y = 16'b0000101100010000;
         4: y = 16'b0000111010111011;
         5: y = 16'b0001001001100011;
         6: y = 16'b0001011000000110;
         7: y = 16'b0001100110100011;
         8: y = 16'b0001110100111001;
         9: y = 16'b0010000011000111;
        10: y = 16'b0010010001001101;
        11: y = 16'b0010011111001010;
        12: y = 16'b0010101100111011;
        13: y = 16'b0010111010100010;
        14: y = 16'b0011000111111100;
        15: y = 16'b0011010101001001;
        16: y = 16'b0011100010001000;
        17: y = 16'b0011101110111000;
        18: y = 16'b0011111011011001;
        19: y = 16'b0100000111101001;
        20: y = 16'b0100010011100111;
        21: y = 16'b0100011111010100;
        22: y = 16'b0100101010101110;
        23: y = 16'b0100110101110011;
        24: y = 16'b0101000000100101;
        25: y = 16'b0101001011000010;
        26: y = 16'b0101010101001000;
        27: y = 16'b0101011110111001;
        28: y = 16'b0101101000010010;
        29: y = 16'b0101110001010011;
        30: y = 16'b0101111001111101;
        31: y = 16'b0110000010001101;
        32: y = 16'b0110001010000100;
        33: y = 16'b0110010001100001;
        34: y = 16'b0110011000100100;
        35: y = 16'b0110011111001011;
        36: y = 16'b0110100101011000;
        37: y = 16'b0110101011001001;
        38: y = 16'b0110110000011101;
        39: y = 16'b0110110101010110;
        40: y = 16'b0110111001110001;
        41: y = 16'b0110111101101111;
        42: y = 16'b0111000001010001;
        43: y = 16'b0111000100010100;
        44: y = 16'b0111000110111010;
        45: y = 16'b0111001001000010;
        46: y = 16'b0111001010101100;
        47: y = 16'b0111001011110111;
        48: y = 16'b0111001100100101;
        49: y = 16'b0111001100110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=349.23Hz, Fs=64453Hz, 16-bit, Volume 100%

module table_64453_F
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 46;

    always_comb
        case (x)
         0: y = 16'b0000000000000000;
         1: y = 16'b0000001111101111;
         2: y = 16'b0000011111011101;
         3: y = 16'b0000101111001000;
         4: y = 16'b0000111110110000;
         5: y = 16'b0001001110010011;
         6: y = 16'b0001011101110000;
         7: y = 16'b0001101101000111;
         8: y = 16'b0001111100010101;
         9: y = 16'b0010001011011010;
        10: y = 16'b0010011010010100;
        11: y = 16'b0010101001000011;
        12: y = 16'b0010110111100110;
        13: y = 16'b0011000101111010;
        14: y = 16'b0011010100000000;
        15: y = 16'b0011100001110110;
        16: y = 16'b0011101111011100;
        17: y = 16'b0011111100101111;
        18: y = 16'b0100001001101111;
        19: y = 16'b0100010110011100;
        20: y = 16'b0100100010110100;
        21: y = 16'b0100101110110110;
        22: y = 16'b0100111010100010;
        23: y = 16'b0101000101110110;
        24: y = 16'b0101010000110010;
        25: y = 16'b0101011011010101;
        26: y = 16'b0101100101011101;
        27: y = 16'b0101101111001011;
        28: y = 16'b0101111000011110;
        29: y = 16'b0110000001010101;
        30: y = 16'b0110001001101111;
        31: y = 16'b0110010001101011;
        32: y = 16'b0110011001001010;
        33: y = 16'b0110100000001001;
        34: y = 16'b0110100110101010;
        35: y = 16'b0110101100101100;
        36: y = 16'b0110110010001101;
        37: y = 16'b0110110111001110;
        38: y = 16'b0110111011101110;
        39: y = 16'b0110111111101101;
        40: y = 16'b0111000011001011;
        41: y = 16'b0111000110000111;
        42: y = 16'b0111001000100001;
        43: y = 16'b0111001010011001;
        44: y = 16'b0111001011101111;
        45: y = 16'b0111001100100011;
        46: y = 16'b0111001100110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=369.99Hz, Fs=64453Hz, 16-bit, Volume 100%

module table_64453_Fs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 44;

    always_comb
        case (x)
         0: y = 16'b0000000000000000;
         1: y = 16'b0000010000011101;
         2: y = 16'b0000100000111000;
         3: y = 16'b0000110001010001;
         4: y = 16'b0001000001100101;
         5: y = 16'b0001010001110100;
         6: y = 16'b0001100001111101;
         7: y = 16'b0001110001111110;
         8: y = 16'b0010000001110101;
         9: y = 16'b0010010001100010;
        10: y = 16'b0010100001000010;
        11: y = 16'b0010110000010110;
        12: y = 16'b0010111111011011;
        13: y = 16'b0011001110010001;
        14: y = 16'b0011011100110110;
        15: y = 16'b0011101011001001;
        16: y = 16'b0011111001001001;
        17: y = 16'b0100000110110100;
        18: y = 16'b0100010100001010;
        19: y = 16'b0100100001001001;
        20: y = 16'b0100101101110001;
        21: y = 16'b0100111010000000;
        22: y = 16'b0101000101110110;
        23: y = 16'b0101010001010001;
        24: y = 16'b0101011100010001;
        25: y = 16'b0101100110110100;
        26: y = 16'b0101110000111010;
        27: y = 16'b0101111010100001;
        28: y = 16'b0110000011101010;
        29: y = 16'b0110001100010100;
        30: y = 16'b0110010100011101;
        31: y = 16'b0110011100000100;
        32: y = 16'b0110100011001011;
        33: y = 16'b0110101001101111;
        34: y = 16'b0110101111110001;
        35: y = 16'b0110110101001111;
        36: y = 16'b0110111010001001;
        37: y = 16'b0110111110100000;
        38: y = 16'b0111000010010010;
        39: y = 16'b0111000101011111;
        40: y = 16'b0111001000001000;
        41: y = 16'b0111001010001011;
        42: y = 16'b0111001011101001;
        43: y = 16'b0111001100100001;
        44: y = 16'b0111001100110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=392.0Hz, Fs=64453Hz, 16-bit, Volume 100%

module table_64453_G
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 41;

    always_comb
        case (x)
         0: y = 16'b0000000000000000;
         1: y = 16'b0000010001101010;
         2: y = 16'b0000100011010010;
         3: y = 16'b0000110100110110;
         4: y = 16'b0001000110010110;
         5: y = 16'b0001010111101111;
         6: y = 16'b0001101001000000;
         7: y = 16'b0001111010000111;
         8: y = 16'b0010001011000010;
         9: y = 16'b0010011011110001;
        10: y = 16'b0010101100010001;
        11: y = 16'b0010111100100000;
        12: y = 16'b0011001100011110;
        13: y = 16'b0011011100001001;
        14: y = 16'b0011101011011111;
        15: y = 16'b0011111010011111;
        16: y = 16'b0100001001000111;
        17: y = 16'b0100010111010111;
        18: y = 16'b0100100101001100;
        19: y = 16'b0100110010100110;
        20: y = 16'b0100111111100011;
        21: y = 16'b0101001100000010;
        22: y = 16'b0101011000000001;
        23: y = 16'b0101100011100001;
        24: y = 16'b0101101110011111;
        25: y = 16'b0101111000111010;
        26: y = 16'b0110000010110011;
        27: y = 16'b0110001100000110;
        28: y = 16'b0110010100110101;
        29: y = 16'b0110011100111110;
        30: y = 16'b0110100100100000;
        31: y = 16'b0110101011011010;
        32: y = 16'b0110110001101100;
        33: y = 16'b0110110111010110;
        34: y = 16'b0110111100010110;
        35: y = 16'b0111000000101100;
        36: y = 16'b0111000100011001;
        37: y = 16'b0111000111011010;
        38: y = 16'b0111001001110001;
        39: y = 16'b0111001011011101;
        40: y = 16'b0111001100011110;
        41: y = 16'b0111001100110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=415.3Hz, Fs=64453Hz, 16-bit, Volume 100%

module table_64453_Gs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 39;

    always_comb
        case (x)
         0: y = 16'b0000000000000000;
         1: y = 16'b0000010010100100;
         2: y = 16'b0000100101000101;
         3: y = 16'b0000110111100011;
         4: y = 16'b0001001001111011;
         5: y = 16'b0001011100001011;
         6: y = 16'b0001101110010010;
         7: y = 16'b0010000000001101;
         8: y = 16'b0010010001111011;
         9: y = 16'b0010100011011010;
        10: y = 16'b0010110100101000;
        11: y = 16'b0011000101100011;
        12: y = 16'b0011010110001010;
        13: y = 16'b0011100110011010;
        14: y = 16'b0011110110010010;
        15: y = 16'b0100000101110001;
        16: y = 16'b0100010100110101;
        17: y = 16'b0100100011011100;
        18: y = 16'b0100110001100101;
        19: y = 16'b0100111111001110;
        20: y = 16'b0101001100010110;
        21: y = 16'b0101011000111011;
        22: y = 16'b0101100100111101;
        23: y = 16'b0101110000011001;
        24: y = 16'b0101111011001111;
        25: y = 16'b0110000101011110;
        26: y = 16'b0110001111000101;
        27: y = 16'b0110011000000010;
        28: y = 16'b0110100000010101;
        29: y = 16'b0110100111111100;
        30: y = 16'b0110101110110111;
        31: y = 16'b0110110101000110;
        32: y = 16'b0110111010101000;
        33: y = 16'b0110111111011011;
        34: y = 16'b0111000011100000;
        35: y = 16'b0111000110110110;
        36: y = 16'b0111001001011101;
        37: y = 16'b0111001011010100;
        38: y = 16'b0111001100011100;
        39: y = 16'b0111001100110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=440.0Hz, Fs=64453Hz, 16-bit, Volume 100%

module table_64453_A
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 37;

    always_comb
        case (x)
         0: y = 16'b0000000000000000;
         1: y = 16'b0000010011100100;
         2: y = 16'b0000100111000101;
         3: y = 16'b0000111010100010;
         4: y = 16'b0001001101111000;
         5: y = 16'b0001100001000101;
         6: y = 16'b0001110100000111;
         7: y = 16'b0010000110111100;
         8: y = 16'b0010011001100001;
         9: y = 16'b0010101011110100;
        10: y = 16'b0010111101110100;
        11: y = 16'b0011001111011101;
        12: y = 16'b0011100000101111;
        13: y = 16'b0011110001100111;
        14: y = 16'b0100000010000011;
        15: y = 16'b0100010010000001;
        16: y = 16'b0100100001011111;
        17: y = 16'b0100110000011101;
        18: y = 16'b0100111110110111;
        19: y = 16'b0101001100101100;
        20: y = 16'b0101011001111011;
        21: y = 16'b0101100110100010;
        22: y = 16'b0101110010011111;
        23: y = 16'b0101111101110010;
        24: y = 16'b0110001000011001;
        25: y = 16'b0110010010010011;
        26: y = 16'b0110011011011110;
        27: y = 16'b0110100011111010;
        28: y = 16'b0110101011100101;
        29: y = 16'b0110110010011111;
        30: y = 16'b0110111000100111;
        31: y = 16'b0110111101111100;
        32: y = 16'b0111000010011110;
        33: y = 16'b0111000110001100;
        34: y = 16'b0111001001000101;
        35: y = 16'b0111001011001010;
        36: y = 16'b0111001100011001;
        37: y = 16'b0111001100110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=466.16Hz, Fs=64453Hz, 16-bit, Volume 100%

module table_64453_As
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 35;

    always_comb
        case (x)
         0: y = 16'b0000000000000000;
         1: y = 16'b0000010100101011;
         2: y = 16'b0000101001010100;
         3: y = 16'b0000111101110111;
         4: y = 16'b0001010010010010;
         5: y = 16'b0001100110100011;
         6: y = 16'b0001111010100110;
         7: y = 16'b0010001110011010;
         8: y = 16'b0010100001111011;
         9: y = 16'b0010110101000111;
        10: y = 16'b0011000111111100;
        11: y = 16'b0011011010010111;
        12: y = 16'b0011101100010110;
        13: y = 16'b0011111101110111;
        14: y = 16'b0100001110110111;
        15: y = 16'b0100011111010100;
        16: y = 16'b0100101111001100;
        17: y = 16'b0100111110011101;
        18: y = 16'b0101001101000101;
        19: y = 16'b0101011011000010;
        20: y = 16'b0101101000010010;
        21: y = 16'b0101110100110100;
        22: y = 16'b0110000000100101;
        23: y = 16'b0110001011100101;
        24: y = 16'b0110010101110011;
        25: y = 16'b0110011111001011;
        26: y = 16'b0110100111101111;
        27: y = 16'b0110101111011011;
        28: y = 16'b0110110110010001;
        29: y = 16'b0110111100001101;
        30: y = 16'b0111000001010001;
        31: y = 16'b0111000101011010;
        32: y = 16'b0111001000101001;
        33: y = 16'b0111001010111101;
        34: y = 16'b0111001100010110;
        35: y = 16'b0111001100110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=493.88Hz, Fs=64453Hz, 16-bit, Volume 100%

module table_64453_B
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 33;

    always_comb
        case (x)
         0: y = 16'b0000000000000000;
         1: y = 16'b0000010101111011;
         2: y = 16'b0000101011110011;
         3: y = 16'b0001000001100101;
         4: y = 16'b0001010111001101;
         5: y = 16'b0001101100101001;
         6: y = 16'b0010000001110101;
         7: y = 16'b0010010110101110;
         8: y = 16'b0010101011010001;
         9: y = 16'b0010111111011011;
        10: y = 16'b0011010011001010;
        11: y = 16'b0011100110011010;
        12: y = 16'b0011111001001001;
        13: y = 16'b0100001011010011;
        14: y = 16'b0100011100110111;
        15: y = 16'b0100101101110001;
        16: y = 16'b0100111110000000;
        17: y = 16'b0101001101100000;
        18: y = 16'b0101011100010001;
        19: y = 16'b0101101010001110;
        20: y = 16'b0101110111010111;
        21: y = 16'b0110000011101010;
        22: y = 16'b0110001111000101;
        23: y = 16'b0110011001100110;
        24: y = 16'b0110100011001011;
        25: y = 16'b0110101011110011;
        26: y = 16'b0110110011011110;
        27: y = 16'b0110111010001001;
        28: y = 16'b0110111111110101;
        29: y = 16'b0111000100011111;
        30: y = 16'b0111001000001000;
        31: y = 16'b0111001010101110;
        32: y = 16'b0111001100010011;
        33: y = 16'b0111001100110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=261.63Hz, Fs=52734Hz, 16-bit, Volume 100%

module table_52734_C
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 50;

    always_comb
        case (x)
         0: y = 16'b0000000000000000;
         1: y = 16'b0000001110011110;
         2: y = 16'b0000011100111100;
         3: y = 16'b0000101011010111;
         4: y = 16'b0000111001110000;
         5: y = 16'b0001001000000110;
         6: y = 16'b0001010110010110;
         7: y = 16'b0001100100100001;
         8: y = 16'b0001110010100110;
         9: y = 16'b0010000000100100;
        10: y = 16'b0010001110011010;
        11: y = 16'b0010011100000110;
        12: y = 16'b0010101001101001;
        13: y = 16'b0010110111000001;
        14: y = 16'b0011000100001101;
        15: y = 16'b0011010001001101;
        16: y = 16'b0011011110000000;
        17: y = 16'b0011101010100101;
        18: y = 16'b0011110110111011;
        19: y = 16'b0100000011000001;
        20: y = 16'b0100001110110111;
        21: y = 16'b0100011010011100;
        22: y = 16'b0100100101101111;
        23: y = 16'b0100110000101111;
        24: y = 16'b0100111011011101;
        25: y = 16'b0101000101110110;
        26: y = 16'b0101001111111011;
        27: y = 16'b0101011001101010;
        28: y = 16'b0101100011000100;
        29: y = 16'b0101101100000111;
        30: y = 16'b0101110100110100;
        31: y = 16'b0101111101001000;
        32: y = 16'b0110000101000101;
        33: y = 16'b0110001100101001;
        34: y = 16'b0110010011110100;
        35: y = 16'b0110011010100110;
        36: y = 16'b0110100000111101;
        37: y = 16'b0110100110111010;
        38: y = 16'b0110101100011101;
        39: y = 16'b0110110001100100;
        40: y = 16'b0110110110010001;
        41: y = 16'b0110111010100001;
        42: y = 16'b0110111110010101;
        43: y = 16'b0111000001101110;
        44: y = 16'b0111000100101010;
        45: y = 16'b0111000111001001;
        46: y = 16'b0111001001001011;
        47: y = 16'b0111001010110001;
        48: y = 16'b0111001011111010;
        49: y = 16'b0111001100100101;
        50: y = 16'b0111001100110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=277.18Hz, Fs=52734Hz, 16-bit, Volume 100%

module table_52734_Cs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 48;

    always_comb
        case (x)
         0: y = 16'b0000000000000000;
         1: y = 16'b0000001111000101;
         2: y = 16'b0000011110001001;
         3: y = 16'b0000101101001011;
         4: y = 16'b0000111100001001;
         5: y = 16'b0001001011000100;
         6: y = 16'b0001011001111010;
         7: y = 16'b0001101000101001;
         8: y = 16'b0001110111010001;
         9: y = 16'b0010000101110001;
        10: y = 16'b0010010100001000;
        11: y = 16'b0010100010010101;
        12: y = 16'b0010110000010110;
        13: y = 16'b0010111110001100;
        14: y = 16'b0011001011110100;
        15: y = 16'b0011011001001110;
        16: y = 16'b0011100110011010;
        17: y = 16'b0011110011010110;
        18: y = 16'b0100000000000001;
        19: y = 16'b0100001100011010;
        20: y = 16'b0100011000100010;
        21: y = 16'b0100100100010110;
        22: y = 16'b0100101111110101;
        23: y = 16'b0100111011000001;
        24: y = 16'b0101000101110110;
        25: y = 16'b0101010000010101;
        26: y = 16'b0101011010011101;
        27: y = 16'b0101100100001110;
        28: y = 16'b0101101101100110;
        29: y = 16'b0101110110100100;
        30: y = 16'b0101111111001010;
        31: y = 16'b0110000111010101;
        32: y = 16'b0110001111000101;
        33: y = 16'b0110010110011010;
        34: y = 16'b0110011101010011;
        35: y = 16'b0110100011101111;
        36: y = 16'b0110101001101111;
        37: y = 16'b0110101111010010;
        38: y = 16'b0110110100010111;
        39: y = 16'b0110111000111110;
        40: y = 16'b0110111101000111;
        41: y = 16'b0111000000110010;
        42: y = 16'b0111000011111101;
        43: y = 16'b0111000110101010;
        44: y = 16'b0111001000111000;
        45: y = 16'b0111001010100110;
        46: y = 16'b0111001011110101;
        47: y = 16'b0111001100100100;
        48: y = 16'b0111001100110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=293.66Hz, Fs=52734Hz, 16-bit, Volume 100%

module table_52734_D
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 45;

    always_comb
        case (x)
         0: y = 16'b0000000000000000;
         1: y = 16'b0000010000000101;
         2: y = 16'b0000100000001001;
         3: y = 16'b0000110000001011;
         4: y = 16'b0001000000001000;
         5: y = 16'b0001010000000001;
         6: y = 16'b0001011111110100;
         7: y = 16'b0001101111011111;
         8: y = 16'b0001111111000001;
         9: y = 16'b0010001110011010;
        10: y = 16'b0010011101100111;
        11: y = 16'b0010101100101000;
        12: y = 16'b0010111011011011;
        13: y = 16'b0011001010000000;
        14: y = 16'b0011011000010110;
        15: y = 16'b0011100110011010;
        16: y = 16'b0011110100001100;
        17: y = 16'b0100000001101100;
        18: y = 16'b0100001110110111;
        19: y = 16'b0100011011101101;
        20: y = 16'b0100101000001101;
        21: y = 16'b0100110100010110;
        22: y = 16'b0101000000000111;
        23: y = 16'b0101001011011111;
        24: y = 16'b0101010110011101;
        25: y = 16'b0101100001000000;
        26: y = 16'b0101101011001000;
        27: y = 16'b0101110100110100;
        28: y = 16'b0101111110000010;
        29: y = 16'b0110000110110011;
        30: y = 16'b0110001111000101;
        31: y = 16'b0110010110111000;
        32: y = 16'b0110011110001011;
        33: y = 16'b0110100100111110;
        34: y = 16'b0110101011010001;
        35: y = 16'b0110110001000001;
        36: y = 16'b0110110110010001;
        37: y = 16'b0110111010111110;
        38: y = 16'b0110111111001000;
        39: y = 16'b0111000010110000;
        40: y = 16'b0111000101110100;
        41: y = 16'b0111001000010101;
        42: y = 16'b0111001010010010;
        43: y = 16'b0111001011101100;
        44: y = 16'b0111001100100010;
        45: y = 16'b0111001100110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=311.13Hz, Fs=52734Hz, 16-bit, Volume 100%

module table_52734_Ds
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 42;

    always_comb
        case (x)
         0: y = 16'b0000000000000000;
         1: y = 16'b0000010001001111;
         2: y = 16'b0000100010011100;
         3: y = 16'b0000110011100110;
         4: y = 16'b0001000100101100;
         5: y = 16'b0001010101101011;
         6: y = 16'b0001100110100011;
         7: y = 16'b0001110111010001;
         8: y = 16'b0010000111110101;
         9: y = 16'b0010011000001101;
        10: y = 16'b0010101000010111;
        11: y = 16'b0010111000010010;
        12: y = 16'b0011000111111100;
        13: y = 16'b0011010111010101;
        14: y = 16'b0011100110011010;
        15: y = 16'b0011110101001011;
        16: y = 16'b0100000011100101;
        17: y = 16'b0100010001101001;
        18: y = 16'b0100011111010100;
        19: y = 16'b0100101100100101;
        20: y = 16'b0100111001011100;
        21: y = 16'b0101000101110110;
        22: y = 16'b0101010001110011;
        23: y = 16'b0101011101010010;
        24: y = 16'b0101101000010010;
        25: y = 16'b0101110010110001;
        26: y = 16'b0101111100101111;
        27: y = 16'b0110000110001100;
        28: y = 16'b0110001111000101;
        29: y = 16'b0110010111011010;
        30: y = 16'b0110011111001011;
        31: y = 16'b0110100110010111;
        32: y = 16'b0110101100111101;
        33: y = 16'b0110110010111101;
        34: y = 16'b0110111000010110;
        35: y = 16'b0110111101000111;
        36: y = 16'b0111000001010001;
        37: y = 16'b0111000100110010;
        38: y = 16'b0111000111101011;
        39: y = 16'b0111001001111011;
        40: y = 16'b0111001011100010;
        41: y = 16'b0111001100011111;
        42: y = 16'b0111001100110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=329.63Hz, Fs=52734Hz, 16-bit, Volume 100%

module table_52734_E
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 40;

    always_comb
        case (x)
         0: y = 16'b0000000000000000;
         1: y = 16'b0000010010000110;
         2: y = 16'b0000100100001010;
         3: y = 16'b0000110110001010;
         4: y = 16'b0001001000000110;
         5: y = 16'b0001011001111010;
         6: y = 16'b0001101011100101;
         7: y = 16'b0001111101000101;
         8: y = 16'b0010001110011010;
         9: y = 16'b0010011111100000;
        10: y = 16'b0010110000010110;
        11: y = 16'b0011000000111011;
        12: y = 16'b0011010001001101;
        13: y = 16'b0011100001001010;
        14: y = 16'b0011110000110010;
        15: y = 16'b0100000000000001;
        16: y = 16'b0100001110110111;
        17: y = 16'b0100011101010010;
        18: y = 16'b0100101011010010;
        19: y = 16'b0100111000110011;
        20: y = 16'b0101000101110110;
        21: y = 16'b0101010010011001;
        22: y = 16'b0101011110011010;
        23: y = 16'b0101101001111001;
        24: y = 16'b0101110100110100;
        25: y = 16'b0101111111001010;
        26: y = 16'b0110001000111010;
        27: y = 16'b0110010010000100;
        28: y = 16'b0110011010100110;
        29: y = 16'b0110100010011111;
        30: y = 16'b0110101001101111;
        31: y = 16'b0110110000010101;
        32: y = 16'b0110110110010001;
        33: y = 16'b0110111011100001;
        34: y = 16'b0111000000000101;
        35: y = 16'b0111000011111101;
        36: y = 16'b0111000111001001;
        37: y = 16'b0111001001101000;
        38: y = 16'b0111001011011001;
        39: y = 16'b0111001100011101;
        40: y = 16'b0111001100110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=349.23Hz, Fs=52734Hz, 16-bit, Volume 100%

module table_52734_F
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 38;

    always_comb
        case (x)
         0: y = 16'b0000000000000000;
         1: y = 16'b0000010011000011;
         2: y = 16'b0000100110000011;
         3: y = 16'b0000111001000000;
         4: y = 16'b0001001011110110;
         5: y = 16'b0001011110100100;
         6: y = 16'b0001110001001000;
         7: y = 16'b0010000011011111;
         8: y = 16'b0010010101101000;
         9: y = 16'b0010100111100001;
        10: y = 16'b0010111001000111;
        11: y = 16'b0011001010011001;
        12: y = 16'b0011011011010101;
        13: y = 16'b0011101011111001;
        14: y = 16'b0011111100000011;
        15: y = 16'b0100001011110001;
        16: y = 16'b0100011011000010;
        17: y = 16'b0100101001110101;
        18: y = 16'b0100111000000110;
        19: y = 16'b0101000101110110;
        20: y = 16'b0101010011000010;
        21: y = 16'b0101011111101001;
        22: y = 16'b0101101011101001;
        23: y = 16'b0101110111000010;
        24: y = 16'b0110000001110010;
        25: y = 16'b0110001011110111;
        26: y = 16'b0110010101010001;
        27: y = 16'b0110011101111111;
        28: y = 16'b0110100110000000;
        29: y = 16'b0110101101010010;
        30: y = 16'b0110110011110110;
        31: y = 16'b0110111001101010;
        32: y = 16'b0110111110101110;
        33: y = 16'b0111000011000000;
        34: y = 16'b0111000110100010;
        35: y = 16'b0111001001010010;
        36: y = 16'b0111001011001111;
        37: y = 16'b0111001100011011;
        38: y = 16'b0111001100110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=369.99Hz, Fs=52734Hz, 16-bit, Volume 100%

module table_52734_Fs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 36;

    always_comb
        case (x)
         0: y = 16'b0000000000000000;
         1: y = 16'b0000010100000110;
         2: y = 16'b0000101000001010;
         3: y = 16'b0000111100001001;
         4: y = 16'b0001010000000001;
         5: y = 16'b0001100011101111;
         6: y = 16'b0001110111010001;
         7: y = 16'b0010001010100100;
         8: y = 16'b0010011101100111;
         9: y = 16'b0010110000010110;
        10: y = 16'b0011000010110000;
        11: y = 16'b0011010100110010;
        12: y = 16'b0011100110011010;
        13: y = 16'b0011110111100110;
        14: y = 16'b0100001000010100;
        15: y = 16'b0100011000100010;
        16: y = 16'b0100101000001101;
        17: y = 16'b0100110111010101;
        18: y = 16'b0101000101110110;
        19: y = 16'b0101010011110000;
        20: y = 16'b0101100001000000;
        21: y = 16'b0101101101100110;
        22: y = 16'b0101111001011110;
        23: y = 16'b0110000100101001;
        24: y = 16'b0110001111000101;
        25: y = 16'b0110011000110000;
        26: y = 16'b0110100001101001;
        27: y = 16'b0110101001101111;
        28: y = 16'b0110110001000001;
        29: y = 16'b0110110111011111;
        30: y = 16'b0110111101000111;
        31: y = 16'b0111000001111001;
        32: y = 16'b0111000101110100;
        33: y = 16'b0111001000111000;
        34: y = 16'b0111001011000100;
        35: y = 16'b0111001100011000;
        36: y = 16'b0111001100110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=392.0Hz, Fs=52734Hz, 16-bit, Volume 100%

module table_52734_G
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 34;

    always_comb
        case (x)
         0: y = 16'b0000000000000000;
         1: y = 16'b0000010101010010;
         2: y = 16'b0000101010100001;
         3: y = 16'b0000111111101011;
         4: y = 16'b0001010100101011;
         5: y = 16'b0001101001100000;
         6: y = 16'b0001111110000111;
         7: y = 16'b0010010010011100;
         8: y = 16'b0010100110011110;
         9: y = 16'b0010111010001000;
        10: y = 16'b0011001101011010;
        11: y = 16'b0011100000001111;
        12: y = 16'b0011110010100110;
        13: y = 16'b0100000100011011;
        14: y = 16'b0100010101101101;
        15: y = 16'b0100100110011001;
        16: y = 16'b0100110110011101;
        17: y = 16'b0101000101110110;
        18: y = 16'b0101010100100011;
        19: y = 16'b0101100010100001;
        20: y = 16'b0101101111101111;
        21: y = 16'b0101111100001011;
        22: y = 16'b0110000111110011;
        23: y = 16'b0110010010100101;
        24: y = 16'b0110011100100000;
        25: y = 16'b0110100101100011;
        26: y = 16'b0110101101101100;
        27: y = 16'b0110110100111011;
        28: y = 16'b0110111011001110;
        29: y = 16'b0111000000100101;
        30: y = 16'b0111000100111110;
        31: y = 16'b0111001000011001;
        32: y = 16'b0111001010110110;
        33: y = 16'b0111001100010101;
        34: y = 16'b0111001100110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=415.3Hz, Fs=52734Hz, 16-bit, Volume 100%

module table_52734_Gs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 32;

    always_comb
        case (x)
         0: y = 16'b0000000000000000;
         1: y = 16'b0000010110100111;
         2: y = 16'b0000101101001011;
         3: y = 16'b0001000011100111;
         4: y = 16'b0001011001111010;
         5: y = 16'b0001101111111110;
         6: y = 16'b0010000101110001;
         7: y = 16'b0010011011010000;
         8: y = 16'b0010110000010110;
         9: y = 16'b0011000101000001;
        10: y = 16'b0011011001001110;
        11: y = 16'b0011101100111010;
        12: y = 16'b0100000000000001;
        13: y = 16'b0100010010100000;
        14: y = 16'b0100100100010110;
        15: y = 16'b0100110101011110;
        16: y = 16'b0101000101110110;
        17: y = 16'b0101010101011100;
        18: y = 16'b0101100100001110;
        19: y = 16'b0101110010001000;
        20: y = 16'b0101111111001010;
        21: y = 16'b0110001011010000;
        22: y = 16'b0110010110011010;
        23: y = 16'b0110100000100100;
        24: y = 16'b0110101001101111;
        25: y = 16'b0110110001111000;
        26: y = 16'b0110111000111110;
        27: y = 16'b0110111111000000;
        28: y = 16'b0111000011111101;
        29: y = 16'b0111000111110101;
        30: y = 16'b0111001010100110;
        31: y = 16'b0111001100010000;
        32: y = 16'b0111001100110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=440.0Hz, Fs=52734Hz, 16-bit, Volume 100%

module table_52734_A
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 30;

    always_comb
        case (x)
         0: y = 16'b0000000000000000;
         1: y = 16'b0000011000000111;
         2: y = 16'b0000110000001011;
         3: y = 16'b0001001000000110;
         4: y = 16'b0001011111110100;
         5: y = 16'b0001110111010001;
         6: y = 16'b0010001110011010;
         7: y = 16'b0010100101001001;
         8: y = 16'b0010111011011011;
         9: y = 16'b0011010001001101;
        10: y = 16'b0011100110011010;
        11: y = 16'b0011111010111110;
        12: y = 16'b0100001110110111;
        13: y = 16'b0100100010000000;
        14: y = 16'b0100110100010110;
        15: y = 16'b0101000101110110;
        16: y = 16'b0101010110011101;
        17: y = 16'b0101100110001000;
        18: y = 16'b0101110100110100;
        19: y = 16'b0110000010011110;
        20: y = 16'b0110001111000101;
        21: y = 16'b0110011010100110;
        22: y = 16'b0110100100111110;
        23: y = 16'b0110101110001101;
        24: y = 16'b0110110110010001;
        25: y = 16'b0110111101000111;
        26: y = 16'b0111000010110000;
        27: y = 16'b0111000111001001;
        28: y = 16'b0111001010010010;
        29: y = 16'b0111001100001100;
        30: y = 16'b0111001100110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=466.16Hz, Fs=52734Hz, 16-bit, Volume 100%

module table_52734_As
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 28;

    always_comb
        case (x)
         0: y = 16'b0000000000000000;
         1: y = 16'b0000011001110110;
         2: y = 16'b0000110011100110;
         3: y = 16'b0001001101001100;
         4: y = 16'b0001100110100011;
         5: y = 16'b0001111111100100;
         6: y = 16'b0010011000001101;
         7: y = 16'b0010110000010110;
         8: y = 16'b0011000111111100;
         9: y = 16'b0011011110111010;
        10: y = 16'b0011110101001011;
        11: y = 16'b0100001010101010;
        12: y = 16'b0100011111010100;
        13: y = 16'b0100110011000100;
        14: y = 16'b0101000101110110;
        15: y = 16'b0101010111100110;
        16: y = 16'b0101101000010010;
        17: y = 16'b0101110111110101;
        18: y = 16'b0110000110001100;
        19: y = 16'b0110010011010100;
        20: y = 16'b0110011111001011;
        21: y = 16'b0110101001101111;
        22: y = 16'b0110110010111101;
        23: y = 16'b0110111010110011;
        24: y = 16'b0111000001010001;
        25: y = 16'b0111000110010011;
        26: y = 16'b0111001001111011;
        27: y = 16'b0111001100000110;
        28: y = 16'b0111001100110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=493.88Hz, Fs=52734Hz, 16-bit, Volume 100%

module table_52734_B
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 27;

    always_comb
        case (x)
         0: y = 16'b0000000000000000;
         1: y = 16'b0000011010110011;
         2: y = 16'b0000110101100000;
         3: y = 16'b0001010000000001;
         4: y = 16'b0001101010010001;
         5: y = 16'b0010000100001010;
         6: y = 16'b0010011101100111;
         7: y = 16'b0010110110100001;
         8: y = 16'b0011001110110100;
         9: y = 16'b0011100110011010;
        10: y = 16'b0011111101001110;
        11: y = 16'b0100010011001011;
        12: y = 16'b0100101000001101;
        13: y = 16'b0100111100001111;
        14: y = 16'b0101001111001100;
        15: y = 16'b0101100001000000;
        16: y = 16'b0101110001101000;
        17: y = 16'b0110000001000000;
        18: y = 16'b0110001111000101;
        19: y = 16'b0110011011110011;
        20: y = 16'b0110100111001000;
        21: y = 16'b0110110001000001;
        22: y = 16'b0110111001011101;
        23: y = 16'b0111000000011001;
        24: y = 16'b0111000101110100;
        25: y = 16'b0111001001101101;
        26: y = 16'b0111001100000010;
        27: y = 16'b0111001100110100;
        default: y = 16'b0;
        endcase

endmodule

