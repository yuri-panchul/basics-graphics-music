`define HUB75E_LED_MATRIX_BRIGHTNESS 8
`include "../tang_primer_25k_pmod_hub75e_led_matrix/board_specific_top.sv"
