// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=261.63Hz, Fs=48828Hz, 16-bit, Volume 15/15 bit

module table_48828_C
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 47;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001111011011;
        2: y = 16'b0000011110110101;
        3: y = 16'b0000101110001101;
        4: y = 16'b0000111101100010;
        5: y = 16'b0001001100110010;
        6: y = 16'b0001011011111101;
        7: y = 16'b0001101011000001;
        8: y = 16'b0001111001111101;
        9: y = 16'b0010001000110001;
        10: y = 16'b0010010111011011;
        11: y = 16'b0010100101111010;
        12: y = 16'b0010110100001110;
        13: y = 16'b0011000010010100;
        14: y = 16'b0011010000001101;
        15: y = 16'b0011011101110110;
        16: y = 16'b0011101011010000;
        17: y = 16'b0011111000011001;
        18: y = 16'b0100000101010000;
        19: y = 16'b0100010001110101;
        20: y = 16'b0100011110000110;
        21: y = 16'b0100101010000010;
        22: y = 16'b0100110101101010;
        23: y = 16'b0101000000111011;
        24: y = 16'b0101001011110101;
        25: y = 16'b0101010110010111;
        26: y = 16'b0101100000100001;
        27: y = 16'b0101101010010010;
        28: y = 16'b0101110011101001;
        29: y = 16'b0101111100100101;
        30: y = 16'b0110000101000110;
        31: y = 16'b0110001101001100;
        32: y = 16'b0110010100110101;
        33: y = 16'b0110011100000001;
        34: y = 16'b0110100010101111;
        35: y = 16'b0110101001000000;
        36: y = 16'b0110101110110010;
        37: y = 16'b0110110100000101;
        38: y = 16'b0110111000111010;
        39: y = 16'b0110111101001110;
        40: y = 16'b0111000001000011;
        41: y = 16'b0111000100011000;
        42: y = 16'b0111000111001100;
        43: y = 16'b0111001001100000;
        44: y = 16'b0111001011010100;
        45: y = 16'b0111001100100110;
        46: y = 16'b0111001101011000;
        47: y = 16'b0111001101101000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=277.18Hz, Fs=48828Hz, 16-bit, Volume 15/15 bit

module table_48828_Cs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 44;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000010000011110;
        2: y = 16'b0000100000111100;
        3: y = 16'b0000110001010110;
        4: y = 16'b0001000001101101;
        5: y = 16'b0001010001111110;
        6: y = 16'b0001100010001000;
        7: y = 16'b0001110010001010;
        8: y = 16'b0010000010000100;
        9: y = 16'b0010010001110010;
        10: y = 16'b0010100001010101;
        11: y = 16'b0010110000101010;
        12: y = 16'b0010111111110001;
        13: y = 16'b0011001110101000;
        14: y = 16'b0011011101001111;
        15: y = 16'b0011101011100011;
        16: y = 16'b0011111001100101;
        17: y = 16'b0100000111010010;
        18: y = 16'b0100010100101001;
        19: y = 16'b0100100001101010;
        20: y = 16'b0100101110010011;
        21: y = 16'b0100111010100100;
        22: y = 16'b0101000110011011;
        23: y = 16'b0101010001110111;
        24: y = 16'b0101011100111000;
        25: y = 16'b0101100111011100;
        26: y = 16'b0101110001100011;
        27: y = 16'b0101111011001100;
        28: y = 16'b0110000100010110;
        29: y = 16'b0110001101000000;
        30: y = 16'b0110010101001010;
        31: y = 16'b0110011100110011;
        32: y = 16'b0110100011111010;
        33: y = 16'b0110101010011111;
        34: y = 16'b0110110000100001;
        35: y = 16'b0110110110000000;
        36: y = 16'b0110111010111011;
        37: y = 16'b0110111111010010;
        38: y = 16'b0111000011000101;
        39: y = 16'b0111000110010011;
        40: y = 16'b0111001000111011;
        41: y = 16'b0111001010111111;
        42: y = 16'b0111001100011101;
        43: y = 16'b0111001101010101;
        44: y = 16'b0111001101101000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=293.66Hz, Fs=48828Hz, 16-bit, Volume 15/15 bit

module table_48828_D
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 42;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000010001010001;
        2: y = 16'b0000100010100000;
        3: y = 16'b0000110011101100;
        4: y = 16'b0001000100110011;
        5: y = 16'b0001010101110101;
        6: y = 16'b0001100110101110;
        7: y = 16'b0001110111011111;
        8: y = 16'b0010001000000100;
        9: y = 16'b0010011000011110;
        10: y = 16'b0010101000101010;
        11: y = 16'b0010111000100110;
        12: y = 16'b0011001000010011;
        13: y = 16'b0011010111101101;
        14: y = 16'b0011100110110100;
        15: y = 16'b0011110101100110;
        16: y = 16'b0100000100000011;
        17: y = 16'b0100010010001000;
        18: y = 16'b0100011111110100;
        19: y = 16'b0100101101000111;
        20: y = 16'b0100111001111111;
        21: y = 16'b0101000110011011;
        22: y = 16'b0101010010011001;
        23: y = 16'b0101011101111010;
        24: y = 16'b0101101000111010;
        25: y = 16'b0101110011011011;
        26: y = 16'b0101111101011010;
        27: y = 16'b0110000110111000;
        28: y = 16'b0110001111110010;
        29: y = 16'b0110011000001000;
        30: y = 16'b0110011111111010;
        31: y = 16'b0110100111000111;
        32: y = 16'b0110101101101110;
        33: y = 16'b0110110011101110;
        34: y = 16'b0110111001000111;
        35: y = 16'b0110111101111001;
        36: y = 16'b0111000010000011;
        37: y = 16'b0111000101100101;
        38: y = 16'b0111001000011110;
        39: y = 16'b0111001010101110;
        40: y = 16'b0111001100010101;
        41: y = 16'b0111001101010011;
        42: y = 16'b0111001101101000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=311.13Hz, Fs=48828Hz, 16-bit, Volume 15/15 bit

module table_48828_Ds
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 39;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000010010100110;
        2: y = 16'b0000100101001001;
        3: y = 16'b0000110111101001;
        4: y = 16'b0001001010000011;
        5: y = 16'b0001011100010110;
        6: y = 16'b0001101110011110;
        7: y = 16'b0010000000011100;
        8: y = 16'b0010010010001100;
        9: y = 16'b0010100011101100;
        10: y = 16'b0010110100111100;
        11: y = 16'b0011000101111001;
        12: y = 16'b0011010110100010;
        13: y = 16'b0011100110110100;
        14: y = 16'b0011110110101110;
        15: y = 16'b0100000110001111;
        16: y = 16'b0100010101010100;
        17: y = 16'b0100100011111101;
        18: y = 16'b0100110010000111;
        19: y = 16'b0100111111110010;
        20: y = 16'b0101001100111011;
        21: y = 16'b0101011001100010;
        22: y = 16'b0101100101100101;
        23: y = 16'b0101110001000011;
        24: y = 16'b0101111011111010;
        25: y = 16'b0110000110001010;
        26: y = 16'b0110001111110010;
        27: y = 16'b0110011000110000;
        28: y = 16'b0110100001000100;
        29: y = 16'b0110101000101100;
        30: y = 16'b0110101111101000;
        31: y = 16'b0110110101111000;
        32: y = 16'b0110111011011010;
        33: y = 16'b0111000000001110;
        34: y = 16'b0111000100010011;
        35: y = 16'b0111000111101001;
        36: y = 16'b0111001010010001;
        37: y = 16'b0111001100001000;
        38: y = 16'b0111001101010000;
        39: y = 16'b0111001101101000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=329.63Hz, Fs=48828Hz, 16-bit, Volume 15/15 bit

module table_48828_E
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 37;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000010011100110;
        2: y = 16'b0000100111001010;
        3: y = 16'b0000111010101001;
        4: y = 16'b0001001110000001;
        5: y = 16'b0001100001010000;
        6: y = 16'b0001110100010100;
        7: y = 16'b0010000111001011;
        8: y = 16'b0010011001110010;
        9: y = 16'b0010101100001000;
        10: y = 16'b0010111110001001;
        11: y = 16'b0011001111110101;
        12: y = 16'b0011100001001000;
        13: y = 16'b0011110010000010;
        14: y = 16'b0100000010100000;
        15: y = 16'b0100010010100000;
        16: y = 16'b0100100010000000;
        17: y = 16'b0100110000111111;
        18: y = 16'b0100111111011011;
        19: y = 16'b0101001101010001;
        20: y = 16'b0101011010100010;
        21: y = 16'b0101100111001010;
        22: y = 16'b0101110011001001;
        23: y = 16'b0101111110011101;
        24: y = 16'b0110001001000110;
        25: y = 16'b0110010011000000;
        26: y = 16'b0110011100001101;
        27: y = 16'b0110100100101001;
        28: y = 16'b0110101100010110;
        29: y = 16'b0110110011010000;
        30: y = 16'b0110111001011001;
        31: y = 16'b0110111110101111;
        32: y = 16'b0111000011010001;
        33: y = 16'b0111000110111111;
        34: y = 16'b0111001001111001;
        35: y = 16'b0111001011111110;
        36: y = 16'b0111001101001101;
        37: y = 16'b0111001101101000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=349.23Hz, Fs=48828Hz, 16-bit, Volume 15/15 bit

module table_48828_F
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 35;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000010100101101;
        2: y = 16'b0000101001011000;
        3: y = 16'b0000111101111110;
        4: y = 16'b0001010010011011;
        5: y = 16'b0001100110101110;
        6: y = 16'b0001111010110100;
        7: y = 16'b0010001110101010;
        8: y = 16'b0010100010001101;
        9: y = 16'b0010110101011100;
        10: y = 16'b0011001000010011;
        11: y = 16'b0011011010110000;
        12: y = 16'b0011101100110001;
        13: y = 16'b0011111110010100;
        14: y = 16'b0100001111010110;
        15: y = 16'b0100011111110100;
        16: y = 16'b0100101111101110;
        17: y = 16'b0100111111000001;
        18: y = 16'b0101001101101010;
        19: y = 16'b0101011011101001;
        20: y = 16'b0101101000111010;
        21: y = 16'b0101110101011110;
        22: y = 16'b0110000001010001;
        23: y = 16'b0110001100010010;
        24: y = 16'b0110010110100000;
        25: y = 16'b0110011111111010;
        26: y = 16'b0110101000011111;
        27: y = 16'b0110110000001100;
        28: y = 16'b0110110111000010;
        29: y = 16'b0110111100111111;
        30: y = 16'b0111000010000011;
        31: y = 16'b0111000110001101;
        32: y = 16'b0111001001011101;
        33: y = 16'b0111001011110001;
        34: y = 16'b0111001101001010;
        35: y = 16'b0111001101101000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=369.99Hz, Fs=48828Hz, 16-bit, Volume 15/15 bit

module table_48828_Fs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 33;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000010101111110;
        2: y = 16'b0000101011111000;
        3: y = 16'b0001000001101101;
        4: y = 16'b0001010111010111;
        5: y = 16'b0001101100110101;
        6: y = 16'b0010000010000100;
        7: y = 16'b0010010110111111;
        8: y = 16'b0010101011100100;
        9: y = 16'b0010111111110001;
        10: y = 16'b0011010011100010;
        11: y = 16'b0011100110110100;
        12: y = 16'b0011111001100101;
        13: y = 16'b0100001011110001;
        14: y = 16'b0100011101010111;
        15: y = 16'b0100101110010011;
        16: y = 16'b0100111110100100;
        17: y = 16'b0101001110000110;
        18: y = 16'b0101011100111000;
        19: y = 16'b0101101010110111;
        20: y = 16'b0101111000000010;
        21: y = 16'b0110000100010110;
        22: y = 16'b0110001111110010;
        23: y = 16'b0110011010010100;
        24: y = 16'b0110100011111010;
        25: y = 16'b0110101100100100;
        26: y = 16'b0110110100001111;
        27: y = 16'b0110111010111011;
        28: y = 16'b0111000000100111;
        29: y = 16'b0111000101010010;
        30: y = 16'b0111001000111011;
        31: y = 16'b0111001011100010;
        32: y = 16'b0111001101000111;
        33: y = 16'b0111001101101000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=392.0Hz, Fs=48828Hz, 16-bit, Volume 15/15 bit

module table_48828_G
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 31;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000010111011000;
        2: y = 16'b0000101110101101;
        3: y = 16'b0001000101111010;
        4: y = 16'b0001011100111011;
        5: y = 16'b0001110011101101;
        6: y = 16'b0010001010001100;
        7: y = 16'b0010100000010101;
        8: y = 16'b0010110110000011;
        9: y = 16'b0011001011010011;
        10: y = 16'b0011100000000010;
        11: y = 16'b0011110100001100;
        12: y = 16'b0100000111101110;
        13: y = 16'b0100011010100100;
        14: y = 16'b0100101100101100;
        15: y = 16'b0100111110000011;
        16: y = 16'b0101001110100101;
        17: y = 16'b0101011110010001;
        18: y = 16'b0101101101000011;
        19: y = 16'b0101111010111001;
        20: y = 16'b0110000111110000;
        21: y = 16'b0110010011101000;
        22: y = 16'b0110011110011101;
        23: y = 16'b0110101000001110;
        24: y = 16'b0110110000111001;
        25: y = 16'b0110111000011101;
        26: y = 16'b0110111110111001;
        27: y = 16'b0111000100001011;
        28: y = 16'b0111001000010011;
        29: y = 16'b0111001011010000;
        30: y = 16'b0111001101000010;
        31: y = 16'b0111001101101000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=415.3Hz, Fs=48828Hz, 16-bit, Volume 15/15 bit

module table_48828_Gs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 29;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000011000111111;
        2: y = 16'b0000110001111010;
        3: y = 16'b0001001010101100;
        4: y = 16'b0001100011001111;
        5: y = 16'b0001111011100000;
        6: y = 16'b0010010011011001;
        7: y = 16'b0010101010110111;
        8: y = 16'b0011000001110101;
        9: y = 16'b0011011000001111;
        10: y = 16'b0011101110000000;
        11: y = 16'b0100000011000100;
        12: y = 16'b0100010111010111;
        13: y = 16'b0100101010110110;
        14: y = 16'b0100111101011101;
        15: y = 16'b0101001111001001;
        16: y = 16'b0101011111110101;
        17: y = 16'b0101101111100000;
        18: y = 16'b0101111110000101;
        19: y = 16'b0110001011100011;
        20: y = 16'b0110010111110110;
        21: y = 16'b0110100010111101;
        22: y = 16'b0110101100110110;
        23: y = 16'b0110110101011101;
        24: y = 16'b0110111100110011;
        25: y = 16'b0111000010110101;
        26: y = 16'b0111000111100011;
        27: y = 16'b0111001010111011;
        28: y = 16'b0111001100111101;
        29: y = 16'b0111001101101000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=440.0Hz, Fs=48828Hz, 16-bit, Volume 15/15 bit

module table_48828_A
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 28;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000011001111001;
        2: y = 16'b0000110011101100;
        3: y = 16'b0001001101010101;
        4: y = 16'b0001100110101110;
        5: y = 16'b0001111111110011;
        6: y = 16'b0010011000011110;
        7: y = 16'b0010110000101010;
        8: y = 16'b0011001000010011;
        9: y = 16'b0011011111010011;
        10: y = 16'b0011110101100110;
        11: y = 16'b0100001011001000;
        12: y = 16'b0100011111110100;
        13: y = 16'b0100110011100111;
        14: y = 16'b0101000110011011;
        15: y = 16'b0101011000001101;
        16: y = 16'b0101101000111010;
        17: y = 16'b0101111000011111;
        18: y = 16'b0110000110111000;
        19: y = 16'b0110010100000010;
        20: y = 16'b0110011111111010;
        21: y = 16'b0110101010011111;
        22: y = 16'b0110110011101110;
        23: y = 16'b0110111011100101;
        24: y = 16'b0111000010000011;
        25: y = 16'b0111000111000111;
        26: y = 16'b0111001010101110;
        27: y = 16'b0111001100111010;
        28: y = 16'b0111001101101000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=466.16Hz, Fs=48828Hz, 16-bit, Volume 15/15 bit

module table_48828_As
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 26;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000011011111000;
        2: y = 16'b0000110111101001;
        3: y = 16'b0001010011001101;
        4: y = 16'b0001101110011110;
        5: y = 16'b0010001001010101;
        6: y = 16'b0010100011101100;
        7: y = 16'b0010111101011101;
        8: y = 16'b0011010110100010;
        9: y = 16'b0011101110110100;
        10: y = 16'b0100000110001111;
        11: y = 16'b0100011100101100;
        12: y = 16'b0100110010000111;
        13: y = 16'b0101000110011011;
        14: y = 16'b0101011001100010;
        15: y = 16'b0101101011011001;
        16: y = 16'b0101111011111010;
        17: y = 16'b0110001011000011;
        18: y = 16'b0110011000110000;
        19: y = 16'b0110100100111101;
        20: y = 16'b0110101111101000;
        21: y = 16'b0110111000101110;
        22: y = 16'b0111000000001110;
        23: y = 16'b0111000110000100;
        24: y = 16'b0111001010010001;
        25: y = 16'b0111001100110010;
        26: y = 16'b0111001101101000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=493.88Hz, Fs=48828Hz, 16-bit, Volume 15/15 bit

module table_48828_B
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 25;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000011100111111;
        2: y = 16'b0000111001110111;
        3: y = 16'b0001010110100000;
        4: y = 16'b0001110010110011;
        5: y = 16'b0010001110101010;
        6: y = 16'b0010101001111100;
        7: y = 16'b0011000100100011;
        8: y = 16'b0011011110011001;
        9: y = 16'b0011110111010110;
        10: y = 16'b0100001111010110;
        11: y = 16'b0100100110010000;
        12: y = 16'b0100111100000000;
        13: y = 16'b0101010000100001;
        14: y = 16'b0101100011101100;
        15: y = 16'b0101110101011110;
        16: y = 16'b0110000101110001;
        17: y = 16'b0110010100100010;
        18: y = 16'b0110100001101100;
        19: y = 16'b0110101101001101;
        20: y = 16'b0110110111000010;
        21: y = 16'b0110111111001000;
        22: y = 16'b0111000101011101;
        23: y = 16'b0111001001111111;
        24: y = 16'b0111001100101110;
        25: y = 16'b0111001101101000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=261.63Hz, Fs=64453Hz, 16-bit, Volume 15/15 bit

module table_64453_C
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 62;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001011101100;
        2: y = 16'b0000010111011000;
        3: y = 16'b0000100011000011;
        4: y = 16'b0000101110101101;
        5: y = 16'b0000111010010101;
        6: y = 16'b0001000101111010;
        7: y = 16'b0001010001011100;
        8: y = 16'b0001011100111011;
        9: y = 16'b0001101000010110;
        10: y = 16'b0001110011101101;
        11: y = 16'b0001111110111111;
        12: y = 16'b0010001010001100;
        13: y = 16'b0010010101010100;
        14: y = 16'b0010100000010101;
        15: y = 16'b0010101011001111;
        16: y = 16'b0010110110000011;
        17: y = 16'b0011000000101111;
        18: y = 16'b0011001011010011;
        19: y = 16'b0011010101101111;
        20: y = 16'b0011100000000010;
        21: y = 16'b0011101010001100;
        22: y = 16'b0011110100001100;
        23: y = 16'b0011111110000010;
        24: y = 16'b0100000111101110;
        25: y = 16'b0100010001001110;
        26: y = 16'b0100011010100100;
        27: y = 16'b0100100011101110;
        28: y = 16'b0100101100101100;
        29: y = 16'b0100110101011110;
        30: y = 16'b0100111110000011;
        31: y = 16'b0101000110011011;
        32: y = 16'b0101001110100101;
        33: y = 16'b0101010110100010;
        34: y = 16'b0101011110010001;
        35: y = 16'b0101100101110001;
        36: y = 16'b0101101101000011;
        37: y = 16'b0101110100000101;
        38: y = 16'b0101111010111001;
        39: y = 16'b0110000001011100;
        40: y = 16'b0110000111110000;
        41: y = 16'b0110001101110100;
        42: y = 16'b0110010011101000;
        43: y = 16'b0110011001001011;
        44: y = 16'b0110011110011101;
        45: y = 16'b0110100011011110;
        46: y = 16'b0110101000001110;
        47: y = 16'b0110101100101100;
        48: y = 16'b0110110000111001;
        49: y = 16'b0110110100110100;
        50: y = 16'b0110111000011101;
        51: y = 16'b0110111011110100;
        52: y = 16'b0110111110111001;
        53: y = 16'b0111000001101011;
        54: y = 16'b0111000100001011;
        55: y = 16'b0111000110011001;
        56: y = 16'b0111001000010011;
        57: y = 16'b0111001001111011;
        58: y = 16'b0111001011010000;
        59: y = 16'b0111001100010011;
        60: y = 16'b0111001101000010;
        61: y = 16'b0111001101011111;
        62: y = 16'b0111001101101000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=277.18Hz, Fs=64453Hz, 16-bit, Volume 15/15 bit

module table_64453_Cs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 58;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001100100000;
        2: y = 16'b0000011000111111;
        3: y = 16'b0000100101011110;
        4: y = 16'b0000110001111010;
        5: y = 16'b0000111110010100;
        6: y = 16'b0001001010101100;
        7: y = 16'b0001010110111111;
        8: y = 16'b0001100011001111;
        9: y = 16'b0001101111011010;
        10: y = 16'b0001111011100000;
        11: y = 16'b0010000111100000;
        12: y = 16'b0010010011011001;
        13: y = 16'b0010011111001100;
        14: y = 16'b0010101010110111;
        15: y = 16'b0010110110011011;
        16: y = 16'b0011000001110101;
        17: y = 16'b0011001101000111;
        18: y = 16'b0011011000001111;
        19: y = 16'b0011100011001100;
        20: y = 16'b0011101110000000;
        21: y = 16'b0011111000100111;
        22: y = 16'b0100000011000100;
        23: y = 16'b0100001101010100;
        24: y = 16'b0100010111010111;
        25: y = 16'b0100100001001110;
        26: y = 16'b0100101010110110;
        27: y = 16'b0100110100010001;
        28: y = 16'b0100111101011101;
        29: y = 16'b0101000110011011;
        30: y = 16'b0101001111001001;
        31: y = 16'b0101010111100111;
        32: y = 16'b0101011111110101;
        33: y = 16'b0101100111110011;
        34: y = 16'b0101101111100000;
        35: y = 16'b0101110110111011;
        36: y = 16'b0101111110000101;
        37: y = 16'b0110000100111101;
        38: y = 16'b0110001011100011;
        39: y = 16'b0110010001110110;
        40: y = 16'b0110010111110110;
        41: y = 16'b0110011101100100;
        42: y = 16'b0110100010111101;
        43: y = 16'b0110101000000100;
        44: y = 16'b0110101100110110;
        45: y = 16'b0110110001010100;
        46: y = 16'b0110110101011101;
        47: y = 16'b0110111001010011;
        48: y = 16'b0110111100110011;
        49: y = 16'b0110111111111111;
        50: y = 16'b0111000010110101;
        51: y = 16'b0111000101010111;
        52: y = 16'b0111000111100011;
        53: y = 16'b0111001001011010;
        54: y = 16'b0111001010111011;
        55: y = 16'b0111001100000111;
        56: y = 16'b0111001100111101;
        57: y = 16'b0111001101011101;
        58: y = 16'b0111001101101000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=293.66Hz, Fs=64453Hz, 16-bit, Volume 15/15 bit

module table_64453_D
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 55;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001101001100;
        2: y = 16'b0000011010010111;
        3: y = 16'b0000100111100000;
        4: y = 16'b0000110100101000;
        5: y = 16'b0001000001101101;
        6: y = 16'b0001001110101110;
        7: y = 16'b0001011011101011;
        8: y = 16'b0001101000100100;
        9: y = 16'b0001110101010111;
        10: y = 16'b0010000010000100;
        11: y = 16'b0010001110101010;
        12: y = 16'b0010011011001000;
        13: y = 16'b0010100111011111;
        14: y = 16'b0010110011101101;
        15: y = 16'b0010111111110001;
        16: y = 16'b0011001011101011;
        17: y = 16'b0011010111011011;
        18: y = 16'b0011100011000000;
        19: y = 16'b0011101110011000;
        20: y = 16'b0011111001100101;
        21: y = 16'b0100000100100100;
        22: y = 16'b0100001111010110;
        23: y = 16'b0100011001111001;
        24: y = 16'b0100100100001110;
        25: y = 16'b0100101110010011;
        26: y = 16'b0100111000001001;
        27: y = 16'b0101000001101110;
        28: y = 16'b0101001011000011;
        29: y = 16'b0101010100000110;
        30: y = 16'b0101011100111000;
        31: y = 16'b0101100101010111;
        32: y = 16'b0101101101100100;
        33: y = 16'b0101110101011110;
        34: y = 16'b0101111101000100;
        35: y = 16'b0110000100010110;
        36: y = 16'b0110001011010100;
        37: y = 16'b0110010001111101;
        38: y = 16'b0110011000010010;
        39: y = 16'b0110011110010001;
        40: y = 16'b0110100011111010;
        41: y = 16'b0110101001001110;
        42: y = 16'b0110101110001011;
        43: y = 16'b0110110010110010;
        44: y = 16'b0110110111000010;
        45: y = 16'b0110111010111011;
        46: y = 16'b0110111110011101;
        47: y = 16'b0111000001101000;
        48: y = 16'b0111000100011100;
        49: y = 16'b0111000110110111;
        50: y = 16'b0111001000111011;
        51: y = 16'b0111001010100111;
        52: y = 16'b0111001011111100;
        53: y = 16'b0111001100111000;
        54: y = 16'b0111001101011100;
        55: y = 16'b0111001101101000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=311.13Hz, Fs=64453Hz, 16-bit, Volume 15/15 bit

module table_64453_Ds
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 52;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001101111100;
        2: y = 16'b0000011011111000;
        3: y = 16'b0000101001110010;
        4: y = 16'b0000110111101001;
        5: y = 16'b0001000101011101;
        6: y = 16'b0001010011001101;
        7: y = 16'b0001100000111001;
        8: y = 16'b0001101110011110;
        9: y = 16'b0001111011111110;
        10: y = 16'b0010001001010101;
        11: y = 16'b0010010110100101;
        12: y = 16'b0010100011101100;
        13: y = 16'b0010110000101010;
        14: y = 16'b0010111101011101;
        15: y = 16'b0011001010000101;
        16: y = 16'b0011010110100010;
        17: y = 16'b0011100010110010;
        18: y = 16'b0011101110110100;
        19: y = 16'b0011111010101001;
        20: y = 16'b0100000110001111;
        21: y = 16'b0100010001100110;
        22: y = 16'b0100011100101100;
        23: y = 16'b0100100111100010;
        24: y = 16'b0100110010000111;
        25: y = 16'b0100111100011010;
        26: y = 16'b0101000110011011;
        27: y = 16'b0101010000001000;
        28: y = 16'b0101011001100010;
        29: y = 16'b0101100010101000;
        30: y = 16'b0101101011011001;
        31: y = 16'b0101110011110100;
        32: y = 16'b0101111011111010;
        33: y = 16'b0110000011101010;
        34: y = 16'b0110001011000011;
        35: y = 16'b0110010010000101;
        36: y = 16'b0110011000110000;
        37: y = 16'b0110011111000011;
        38: y = 16'b0110100100111101;
        39: y = 16'b0110101010011111;
        40: y = 16'b0110101111101000;
        41: y = 16'b0110110100011000;
        42: y = 16'b0110111000101110;
        43: y = 16'b0110111100101011;
        44: y = 16'b0111000000001110;
        45: y = 16'b0111000011010110;
        46: y = 16'b0111000110000100;
        47: y = 16'b0111001000011000;
        48: y = 16'b0111001010010001;
        49: y = 16'b0111001011101111;
        50: y = 16'b0111001100110010;
        51: y = 16'b0111001101011011;
        52: y = 16'b0111001101101000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=329.63Hz, Fs=64453Hz, 16-bit, Volume 15/15 bit

module table_64453_E
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 49;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001110110011;
        2: y = 16'b0000011101100101;
        3: y = 16'b0000101100010101;
        4: y = 16'b0000111011000010;
        5: y = 16'b0001001001101011;
        6: y = 16'b0001011000010000;
        7: y = 16'b0001100110101110;
        8: y = 16'b0001110101000110;
        9: y = 16'b0010000011010110;
        10: y = 16'b0010010001011110;
        11: y = 16'b0010011111011011;
        12: y = 16'b0010101101001111;
        13: y = 16'b0010111010110111;
        14: y = 16'b0011001000010011;
        15: y = 16'b0011010101100001;
        16: y = 16'b0011100010100010;
        17: y = 16'b0011101111010011;
        18: y = 16'b0011111011110101;
        19: y = 16'b0100001000000111;
        20: y = 16'b0100010100000111;
        21: y = 16'b0100011111110100;
        22: y = 16'b0100101011001111;
        23: y = 16'b0100110110010110;
        24: y = 16'b0101000001001001;
        25: y = 16'b0101001011100111;
        26: y = 16'b0101010101101111;
        27: y = 16'b0101011111100000;
        28: y = 16'b0101101000111010;
        29: y = 16'b0101110001111101;
        30: y = 16'b0101111010100111;
        31: y = 16'b0110000010111000;
        32: y = 16'b0110001010110000;
        33: y = 16'b0110010010001110;
        34: y = 16'b0110011001010010;
        35: y = 16'b0110011111111010;
        36: y = 16'b0110100110000111;
        37: y = 16'b0110101011111001;
        38: y = 16'b0110110001001110;
        39: y = 16'b0110110110000111;
        40: y = 16'b0110111010100011;
        41: y = 16'b0110111110100010;
        42: y = 16'b0111000010000011;
        43: y = 16'b0111000101000111;
        44: y = 16'b0111000111101101;
        45: y = 16'b0111001001110101;
        46: y = 16'b0111001011011111;
        47: y = 16'b0111001100101011;
        48: y = 16'b0111001101011001;
        49: y = 16'b0111001101101000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=349.23Hz, Fs=64453Hz, 16-bit, Volume 15/15 bit

module table_64453_F
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 46;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001111110001;
        2: y = 16'b0000011111100000;
        3: y = 16'b0000101111001101;
        4: y = 16'b0000111110110111;
        5: y = 16'b0001001110011100;
        6: y = 16'b0001011101111011;
        7: y = 16'b0001101101010011;
        8: y = 16'b0001111100100011;
        9: y = 16'b0010001011101001;
        10: y = 16'b0010011010100110;
        11: y = 16'b0010101001010110;
        12: y = 16'b0010110111111010;
        13: y = 16'b0011000110010001;
        14: y = 16'b0011010100011000;
        15: y = 16'b0011100010010000;
        16: y = 16'b0011101111110111;
        17: y = 16'b0011111101001011;
        18: y = 16'b0100001010001101;
        19: y = 16'b0100010110111100;
        20: y = 16'b0100100011010101;
        21: y = 16'b0100101111011000;
        22: y = 16'b0100111011000101;
        23: y = 16'b0101000110011011;
        24: y = 16'b0101010001011000;
        25: y = 16'b0101011011111100;
        26: y = 16'b0101100110000110;
        27: y = 16'b0101101111110101;
        28: y = 16'b0101111001001001;
        29: y = 16'b0110000010000000;
        30: y = 16'b0110001010011011;
        31: y = 16'b0110010010011000;
        32: y = 16'b0110011001111000;
        33: y = 16'b0110100000111000;
        34: y = 16'b0110100111011010;
        35: y = 16'b0110101101011100;
        36: y = 16'b0110110010111110;
        37: y = 16'b0110111000000000;
        38: y = 16'b0110111100100000;
        39: y = 16'b0111000000100000;
        40: y = 16'b0111000011111110;
        41: y = 16'b0111000110111010;
        42: y = 16'b0111001001010101;
        43: y = 16'b0111001011001101;
        44: y = 16'b0111001100100011;
        45: y = 16'b0111001101010111;
        46: y = 16'b0111001101101000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=369.99Hz, Fs=64453Hz, 16-bit, Volume 15/15 bit

module table_64453_Fs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 44;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000010000011110;
        2: y = 16'b0000100000111100;
        3: y = 16'b0000110001010110;
        4: y = 16'b0001000001101101;
        5: y = 16'b0001010001111110;
        6: y = 16'b0001100010001000;
        7: y = 16'b0001110010001010;
        8: y = 16'b0010000010000100;
        9: y = 16'b0010010001110010;
        10: y = 16'b0010100001010101;
        11: y = 16'b0010110000101010;
        12: y = 16'b0010111111110001;
        13: y = 16'b0011001110101000;
        14: y = 16'b0011011101001111;
        15: y = 16'b0011101011100011;
        16: y = 16'b0011111001100101;
        17: y = 16'b0100000111010010;
        18: y = 16'b0100010100101001;
        19: y = 16'b0100100001101010;
        20: y = 16'b0100101110010011;
        21: y = 16'b0100111010100100;
        22: y = 16'b0101000110011011;
        23: y = 16'b0101010001110111;
        24: y = 16'b0101011100111000;
        25: y = 16'b0101100111011100;
        26: y = 16'b0101110001100011;
        27: y = 16'b0101111011001100;
        28: y = 16'b0110000100010110;
        29: y = 16'b0110001101000000;
        30: y = 16'b0110010101001010;
        31: y = 16'b0110011100110011;
        32: y = 16'b0110100011111010;
        33: y = 16'b0110101010011111;
        34: y = 16'b0110110000100001;
        35: y = 16'b0110110110000000;
        36: y = 16'b0110111010111011;
        37: y = 16'b0110111111010010;
        38: y = 16'b0111000011000101;
        39: y = 16'b0111000110010011;
        40: y = 16'b0111001000111011;
        41: y = 16'b0111001010111111;
        42: y = 16'b0111001100011101;
        43: y = 16'b0111001101010101;
        44: y = 16'b0111001101101000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=392.0Hz, Fs=64453Hz, 16-bit, Volume 15/15 bit

module table_64453_G
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 41;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000010001101100;
        2: y = 16'b0000100011010110;
        3: y = 16'b0000110100111100;
        4: y = 16'b0001000110011110;
        5: y = 16'b0001010111111001;
        6: y = 16'b0001101001001100;
        7: y = 16'b0001111010010101;
        8: y = 16'b0010001011010010;
        9: y = 16'b0010011100000010;
        10: y = 16'b0010101100100100;
        11: y = 16'b0010111100110110;
        12: y = 16'b0011001100110101;
        13: y = 16'b0011011100100010;
        14: y = 16'b0011101011111010;
        15: y = 16'b0011111010111011;
        16: y = 16'b0100001001100101;
        17: y = 16'b0100010111110110;
        18: y = 16'b0100100101101101;
        19: y = 16'b0100110011001000;
        20: y = 16'b0101000000000111;
        21: y = 16'b0101001100100111;
        22: y = 16'b0101011000101000;
        23: y = 16'b0101100100001001;
        24: y = 16'b0101101111001000;
        25: y = 16'b0101111001100101;
        26: y = 16'b0110000011011110;
        27: y = 16'b0110001100110011;
        28: y = 16'b0110010101100011;
        29: y = 16'b0110011101101100;
        30: y = 16'b0110100101001111;
        31: y = 16'b0110101100001010;
        32: y = 16'b0110110010011101;
        33: y = 16'b0110111000000111;
        34: y = 16'b0110111101001000;
        35: y = 16'b0111000001011111;
        36: y = 16'b0111000101001100;
        37: y = 16'b0111001000001110;
        38: y = 16'b0111001010100101;
        39: y = 16'b0111001100010001;
        40: y = 16'b0111001101010010;
        41: y = 16'b0111001101101000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=415.3Hz, Fs=64453Hz, 16-bit, Volume 15/15 bit

module table_64453_Gs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 39;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000010010100110;
        2: y = 16'b0000100101001001;
        3: y = 16'b0000110111101001;
        4: y = 16'b0001001010000011;
        5: y = 16'b0001011100010110;
        6: y = 16'b0001101110011110;
        7: y = 16'b0010000000011100;
        8: y = 16'b0010010010001100;
        9: y = 16'b0010100011101100;
        10: y = 16'b0010110100111100;
        11: y = 16'b0011000101111001;
        12: y = 16'b0011010110100010;
        13: y = 16'b0011100110110100;
        14: y = 16'b0011110110101110;
        15: y = 16'b0100000110001111;
        16: y = 16'b0100010101010100;
        17: y = 16'b0100100011111101;
        18: y = 16'b0100110010000111;
        19: y = 16'b0100111111110010;
        20: y = 16'b0101001100111011;
        21: y = 16'b0101011001100010;
        22: y = 16'b0101100101100101;
        23: y = 16'b0101110001000011;
        24: y = 16'b0101111011111010;
        25: y = 16'b0110000110001010;
        26: y = 16'b0110001111110010;
        27: y = 16'b0110011000110000;
        28: y = 16'b0110100001000100;
        29: y = 16'b0110101000101100;
        30: y = 16'b0110101111101000;
        31: y = 16'b0110110101111000;
        32: y = 16'b0110111011011010;
        33: y = 16'b0111000000001110;
        34: y = 16'b0111000100010011;
        35: y = 16'b0111000111101001;
        36: y = 16'b0111001010010001;
        37: y = 16'b0111001100001000;
        38: y = 16'b0111001101010000;
        39: y = 16'b0111001101101000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=440.0Hz, Fs=64453Hz, 16-bit, Volume 15/15 bit

module table_64453_A
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 37;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000010011100110;
        2: y = 16'b0000100111001010;
        3: y = 16'b0000111010101001;
        4: y = 16'b0001001110000001;
        5: y = 16'b0001100001010000;
        6: y = 16'b0001110100010100;
        7: y = 16'b0010000111001011;
        8: y = 16'b0010011001110010;
        9: y = 16'b0010101100001000;
        10: y = 16'b0010111110001001;
        11: y = 16'b0011001111110101;
        12: y = 16'b0011100001001000;
        13: y = 16'b0011110010000010;
        14: y = 16'b0100000010100000;
        15: y = 16'b0100010010100000;
        16: y = 16'b0100100010000000;
        17: y = 16'b0100110000111111;
        18: y = 16'b0100111111011011;
        19: y = 16'b0101001101010001;
        20: y = 16'b0101011010100010;
        21: y = 16'b0101100111001010;
        22: y = 16'b0101110011001001;
        23: y = 16'b0101111110011101;
        24: y = 16'b0110001001000110;
        25: y = 16'b0110010011000000;
        26: y = 16'b0110011100001101;
        27: y = 16'b0110100100101001;
        28: y = 16'b0110101100010110;
        29: y = 16'b0110110011010000;
        30: y = 16'b0110111001011001;
        31: y = 16'b0110111110101111;
        32: y = 16'b0111000011010001;
        33: y = 16'b0111000110111111;
        34: y = 16'b0111001001111001;
        35: y = 16'b0111001011111110;
        36: y = 16'b0111001101001101;
        37: y = 16'b0111001101101000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=466.16Hz, Fs=64453Hz, 16-bit, Volume 15/15 bit

module table_64453_As
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 35;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000010100101101;
        2: y = 16'b0000101001011000;
        3: y = 16'b0000111101111110;
        4: y = 16'b0001010010011011;
        5: y = 16'b0001100110101110;
        6: y = 16'b0001111010110100;
        7: y = 16'b0010001110101010;
        8: y = 16'b0010100010001101;
        9: y = 16'b0010110101011100;
        10: y = 16'b0011001000010011;
        11: y = 16'b0011011010110000;
        12: y = 16'b0011101100110001;
        13: y = 16'b0011111110010100;
        14: y = 16'b0100001111010110;
        15: y = 16'b0100011111110100;
        16: y = 16'b0100101111101110;
        17: y = 16'b0100111111000001;
        18: y = 16'b0101001101101010;
        19: y = 16'b0101011011101001;
        20: y = 16'b0101101000111010;
        21: y = 16'b0101110101011110;
        22: y = 16'b0110000001010001;
        23: y = 16'b0110001100010010;
        24: y = 16'b0110010110100000;
        25: y = 16'b0110011111111010;
        26: y = 16'b0110101000011111;
        27: y = 16'b0110110000001100;
        28: y = 16'b0110110111000010;
        29: y = 16'b0110111100111111;
        30: y = 16'b0111000010000011;
        31: y = 16'b0111000110001101;
        32: y = 16'b0111001001011101;
        33: y = 16'b0111001011110001;
        34: y = 16'b0111001101001010;
        35: y = 16'b0111001101101000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=493.88Hz, Fs=64453Hz, 16-bit, Volume 15/15 bit

module table_64453_B
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 33;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000010101111110;
        2: y = 16'b0000101011111000;
        3: y = 16'b0001000001101101;
        4: y = 16'b0001010111010111;
        5: y = 16'b0001101100110101;
        6: y = 16'b0010000010000100;
        7: y = 16'b0010010110111111;
        8: y = 16'b0010101011100100;
        9: y = 16'b0010111111110001;
        10: y = 16'b0011010011100010;
        11: y = 16'b0011100110110100;
        12: y = 16'b0011111001100101;
        13: y = 16'b0100001011110001;
        14: y = 16'b0100011101010111;
        15: y = 16'b0100101110010011;
        16: y = 16'b0100111110100100;
        17: y = 16'b0101001110000110;
        18: y = 16'b0101011100111000;
        19: y = 16'b0101101010110111;
        20: y = 16'b0101111000000010;
        21: y = 16'b0110000100010110;
        22: y = 16'b0110001111110010;
        23: y = 16'b0110011010010100;
        24: y = 16'b0110100011111010;
        25: y = 16'b0110101100100100;
        26: y = 16'b0110110100001111;
        27: y = 16'b0110111010111011;
        28: y = 16'b0111000000100111;
        29: y = 16'b0111000101010010;
        30: y = 16'b0111001000111011;
        31: y = 16'b0111001011100010;
        32: y = 16'b0111001101000111;
        33: y = 16'b0111001101101000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=261.63Hz, Fs=52734Hz, 16-bit, Volume 15/15 bit

module table_52734_C
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 50;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001110100000;
        2: y = 16'b0000011100111111;
        3: y = 16'b0000101011011100;
        4: y = 16'b0000111001110111;
        5: y = 16'b0001001000001110;
        6: y = 16'b0001010110100000;
        7: y = 16'b0001100100101101;
        8: y = 16'b0001110010110011;
        9: y = 16'b0010000000110011;
        10: y = 16'b0010001110101010;
        11: y = 16'b0010011100011000;
        12: y = 16'b0010101001111100;
        13: y = 16'b0010110111010101;
        14: y = 16'b0011000100100011;
        15: y = 16'b0011010001100101;
        16: y = 16'b0011011110011001;
        17: y = 16'b0011101010111111;
        18: y = 16'b0011110111010110;
        19: y = 16'b0100000011011110;
        20: y = 16'b0100001111010110;
        21: y = 16'b0100011010111100;
        22: y = 16'b0100100110010000;
        23: y = 16'b0100110001010010;
        24: y = 16'b0100111100000000;
        25: y = 16'b0101000110011011;
        26: y = 16'b0101010000100001;
        27: y = 16'b0101011010010001;
        28: y = 16'b0101100011101100;
        29: y = 16'b0101101100110000;
        30: y = 16'b0101110101011110;
        31: y = 16'b0101111101110011;
        32: y = 16'b0110000101110001;
        33: y = 16'b0110001101010110;
        34: y = 16'b0110010100100010;
        35: y = 16'b0110011011010100;
        36: y = 16'b0110100001101100;
        37: y = 16'b0110100111101010;
        38: y = 16'b0110101101001101;
        39: y = 16'b0110110010010101;
        40: y = 16'b0110110111000010;
        41: y = 16'b0110111011010011;
        42: y = 16'b0110111111001000;
        43: y = 16'b0111000010100000;
        44: y = 16'b0111000101011101;
        45: y = 16'b0111000111111100;
        46: y = 16'b0111001001111111;
        47: y = 16'b0111001011100101;
        48: y = 16'b0111001100101110;
        49: y = 16'b0111001101011001;
        50: y = 16'b0111001101101000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=277.18Hz, Fs=52734Hz, 16-bit, Volume 15/15 bit

module table_52734_Cs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 48;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001111000111;
        2: y = 16'b0000011110001100;
        3: y = 16'b0000101101010000;
        4: y = 16'b0000111100010000;
        5: y = 16'b0001001011001101;
        6: y = 16'b0001011010000100;
        7: y = 16'b0001101000110101;
        8: y = 16'b0001110111011111;
        9: y = 16'b0010000110000000;
        10: y = 16'b0010010100011001;
        11: y = 16'b0010100010100111;
        12: y = 16'b0010110000101010;
        13: y = 16'b0010111110100001;
        14: y = 16'b0011001100001011;
        15: y = 16'b0011011001100111;
        16: y = 16'b0011100110110100;
        17: y = 16'b0011110011110001;
        18: y = 16'b0100000000011110;
        19: y = 16'b0100001100111001;
        20: y = 16'b0100011001000001;
        21: y = 16'b0100100100110111;
        22: y = 16'b0100110000011000;
        23: y = 16'b0100111011100100;
        24: y = 16'b0101000110011011;
        25: y = 16'b0101010000111011;
        26: y = 16'b0101011011000100;
        27: y = 16'b0101100100110110;
        28: y = 16'b0101101110001111;
        29: y = 16'b0101110111001111;
        30: y = 16'b0101111111110101;
        31: y = 16'b0110001000000001;
        32: y = 16'b0110001111110010;
        33: y = 16'b0110010111000111;
        34: y = 16'b0110011110000001;
        35: y = 16'b0110100100011111;
        36: y = 16'b0110101010011111;
        37: y = 16'b0110110000000010;
        38: y = 16'b0110110101001000;
        39: y = 16'b0110111001110000;
        40: y = 16'b0110111101111001;
        41: y = 16'b0111000001100100;
        42: y = 16'b0111000100110000;
        43: y = 16'b0111000111011101;
        44: y = 16'b0111001001101011;
        45: y = 16'b0111001011011010;
        46: y = 16'b0111001100101001;
        47: y = 16'b0111001101011000;
        48: y = 16'b0111001101101000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=293.66Hz, Fs=52734Hz, 16-bit, Volume 15/15 bit

module table_52734_D
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 45;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000010000000111;
        2: y = 16'b0000100000001101;
        3: y = 16'b0000110000010000;
        4: y = 16'b0001000000010000;
        5: y = 16'b0001010000001010;
        6: y = 16'b0001011111111111;
        7: y = 16'b0001101111101011;
        8: y = 16'b0001111111001111;
        9: y = 16'b0010001110101010;
        10: y = 16'b0010011101111001;
        11: y = 16'b0010101100111011;
        12: y = 16'b0010111011110001;
        13: y = 16'b0011001010010111;
        14: y = 16'b0011011000101110;
        15: y = 16'b0011100110110100;
        16: y = 16'b0011110100101000;
        17: y = 16'b0100000010001001;
        18: y = 16'b0100001111010110;
        19: y = 16'b0100011100001101;
        20: y = 16'b0100101000101111;
        21: y = 16'b0100110100111001;
        22: y = 16'b0101000000101011;
        23: y = 16'b0101001100000100;
        24: y = 16'b0101010111000011;
        25: y = 16'b0101100001101000;
        26: y = 16'b0101101011110001;
        27: y = 16'b0101110101011110;
        28: y = 16'b0101111110101101;
        29: y = 16'b0110000111011111;
        30: y = 16'b0110001111110010;
        31: y = 16'b0110010111100110;
        32: y = 16'b0110011110111010;
        33: y = 16'b0110100101101110;
        34: y = 16'b0110101100000001;
        35: y = 16'b0110110001110010;
        36: y = 16'b0110110111000010;
        37: y = 16'b0110111011110000;
        38: y = 16'b0110111111111010;
        39: y = 16'b0111000011100010;
        40: y = 16'b0111000110100111;
        41: y = 16'b0111001001001000;
        42: y = 16'b0111001011000110;
        43: y = 16'b0111001100100000;
        44: y = 16'b0111001101010110;
        45: y = 16'b0111001101101000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=311.13Hz, Fs=52734Hz, 16-bit, Volume 15/15 bit

module table_52734_Ds
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 42;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000010001010001;
        2: y = 16'b0000100010100000;
        3: y = 16'b0000110011101100;
        4: y = 16'b0001000100110011;
        5: y = 16'b0001010101110101;
        6: y = 16'b0001100110101110;
        7: y = 16'b0001110111011111;
        8: y = 16'b0010001000000100;
        9: y = 16'b0010011000011110;
        10: y = 16'b0010101000101010;
        11: y = 16'b0010111000100110;
        12: y = 16'b0011001000010011;
        13: y = 16'b0011010111101101;
        14: y = 16'b0011100110110100;
        15: y = 16'b0011110101100110;
        16: y = 16'b0100000100000011;
        17: y = 16'b0100010010001000;
        18: y = 16'b0100011111110100;
        19: y = 16'b0100101101000111;
        20: y = 16'b0100111001111111;
        21: y = 16'b0101000110011011;
        22: y = 16'b0101010010011001;
        23: y = 16'b0101011101111010;
        24: y = 16'b0101101000111010;
        25: y = 16'b0101110011011011;
        26: y = 16'b0101111101011010;
        27: y = 16'b0110000110111000;
        28: y = 16'b0110001111110010;
        29: y = 16'b0110011000001000;
        30: y = 16'b0110011111111010;
        31: y = 16'b0110100111000111;
        32: y = 16'b0110101101101110;
        33: y = 16'b0110110011101110;
        34: y = 16'b0110111001000111;
        35: y = 16'b0110111101111001;
        36: y = 16'b0111000010000011;
        37: y = 16'b0111000101100101;
        38: y = 16'b0111001000011110;
        39: y = 16'b0111001010101110;
        40: y = 16'b0111001100010101;
        41: y = 16'b0111001101010011;
        42: y = 16'b0111001101101000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=329.63Hz, Fs=52734Hz, 16-bit, Volume 15/15 bit

module table_52734_E
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 40;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000010010001000;
        2: y = 16'b0000100100001110;
        3: y = 16'b0000110110010001;
        4: y = 16'b0001001000001110;
        5: y = 16'b0001011010000100;
        6: y = 16'b0001101011110001;
        7: y = 16'b0001111101010011;
        8: y = 16'b0010001110101010;
        9: y = 16'b0010011111110010;
        10: y = 16'b0010110000101010;
        11: y = 16'b0011000001010001;
        12: y = 16'b0011010001100101;
        13: y = 16'b0011100001100100;
        14: y = 16'b0011110001001101;
        15: y = 16'b0100000000011110;
        16: y = 16'b0100001111010110;
        17: y = 16'b0100011101110011;
        18: y = 16'b0100101011110011;
        19: y = 16'b0100111001010110;
        20: y = 16'b0101000110011011;
        21: y = 16'b0101010010111111;
        22: y = 16'b0101011111000001;
        23: y = 16'b0101101010100001;
        24: y = 16'b0101110101011110;
        25: y = 16'b0101111111110101;
        26: y = 16'b0110001001100110;
        27: y = 16'b0110010010110001;
        28: y = 16'b0110011011010100;
        29: y = 16'b0110100011001110;
        30: y = 16'b0110101010011111;
        31: y = 16'b0110110001000110;
        32: y = 16'b0110110111000010;
        33: y = 16'b0110111100010011;
        34: y = 16'b0111000000111000;
        35: y = 16'b0111000100110000;
        36: y = 16'b0111000111111100;
        37: y = 16'b0111001010011011;
        38: y = 16'b0111001100001101;
        39: y = 16'b0111001101010001;
        40: y = 16'b0111001101101000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=349.23Hz, Fs=52734Hz, 16-bit, Volume 15/15 bit

module table_52734_F
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 38;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000010011000101;
        2: y = 16'b0000100110001000;
        3: y = 16'b0000111001000110;
        4: y = 16'b0001001011111111;
        5: y = 16'b0001011110101111;
        6: y = 16'b0001110001010101;
        7: y = 16'b0010000011101110;
        8: y = 16'b0010010101111001;
        9: y = 16'b0010100111110011;
        10: y = 16'b0010111001011100;
        11: y = 16'b0011001010110000;
        12: y = 16'b0011011011101101;
        13: y = 16'b0011101100010011;
        14: y = 16'b0011111100011111;
        15: y = 16'b0100001100001111;
        16: y = 16'b0100011011100010;
        17: y = 16'b0100101010010110;
        18: y = 16'b0100111000101010;
        19: y = 16'b0101000110011011;
        20: y = 16'b0101010011101000;
        21: y = 16'b0101100000010001;
        22: y = 16'b0101101100010010;
        23: y = 16'b0101110111101100;
        24: y = 16'b0110000010011101;
        25: y = 16'b0110001100100100;
        26: y = 16'b0110010101111111;
        27: y = 16'b0110011110101110;
        28: y = 16'b0110100110110000;
        29: y = 16'b0110101110000011;
        30: y = 16'b0110110100100111;
        31: y = 16'b0110111010011100;
        32: y = 16'b0110111111100000;
        33: y = 16'b0111000011110011;
        34: y = 16'b0111000111010101;
        35: y = 16'b0111001010000101;
        36: y = 16'b0111001100000011;
        37: y = 16'b0111001101001111;
        38: y = 16'b0111001101101000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=369.99Hz, Fs=52734Hz, 16-bit, Volume 15/15 bit

module table_52734_Fs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 36;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000010100001001;
        2: y = 16'b0000101000001111;
        3: y = 16'b0000111100010000;
        4: y = 16'b0001010000001010;
        5: y = 16'b0001100011111010;
        6: y = 16'b0001110111011111;
        7: y = 16'b0010001010110100;
        8: y = 16'b0010011101111001;
        9: y = 16'b0010110000101010;
        10: y = 16'b0011000011000110;
        11: y = 16'b0011010101001010;
        12: y = 16'b0011100110110100;
        13: y = 16'b0011111000000010;
        14: y = 16'b0100001000110010;
        15: y = 16'b0100011001000001;
        16: y = 16'b0100101000101111;
        17: y = 16'b0100110111111000;
        18: y = 16'b0101000110011011;
        19: y = 16'b0101010100010110;
        20: y = 16'b0101100001101000;
        21: y = 16'b0101101110001111;
        22: y = 16'b0101111010001001;
        23: y = 16'b0110000101010101;
        24: y = 16'b0110001111110010;
        25: y = 16'b0110011001011110;
        26: y = 16'b0110100010011000;
        27: y = 16'b0110101010011111;
        28: y = 16'b0110110001110010;
        29: y = 16'b0110111000010001;
        30: y = 16'b0110111101111001;
        31: y = 16'b0111000010101100;
        32: y = 16'b0111000110100111;
        33: y = 16'b0111001001101011;
        34: y = 16'b0111001011111000;
        35: y = 16'b0111001101001100;
        36: y = 16'b0111001101101000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=392.0Hz, Fs=52734Hz, 16-bit, Volume 15/15 bit

module table_52734_G
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 34;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000010101010100;
        2: y = 16'b0000101010100110;
        3: y = 16'b0000111111110010;
        4: y = 16'b0001010100110101;
        5: y = 16'b0001101001101100;
        6: y = 16'b0001111110010101;
        7: y = 16'b0010010010101101;
        8: y = 16'b0010100110110001;
        9: y = 16'b0010111010011101;
        10: y = 16'b0011001101110001;
        11: y = 16'b0011100000101000;
        12: y = 16'b0011110011000001;
        13: y = 16'b0100000100111000;
        14: y = 16'b0100010110001100;
        15: y = 16'b0100100110111010;
        16: y = 16'b0100110111000000;
        17: y = 16'b0101000110011011;
        18: y = 16'b0101010101001001;
        19: y = 16'b0101100011001001;
        20: y = 16'b0101110000011001;
        21: y = 16'b0101111100110110;
        22: y = 16'b0110001000011111;
        23: y = 16'b0110010011010010;
        24: y = 16'b0110011101001111;
        25: y = 16'b0110100110010011;
        26: y = 16'b0110101110011101;
        27: y = 16'b0110110101101100;
        28: y = 16'b0110111100000000;
        29: y = 16'b0111000001010111;
        30: y = 16'b0111000101110001;
        31: y = 16'b0111001001001101;
        32: y = 16'b0111001011101010;
        33: y = 16'b0111001101001000;
        34: y = 16'b0111001101101000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=415.3Hz, Fs=52734Hz, 16-bit, Volume 15/15 bit

module table_52734_Gs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 32;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000010110101010;
        2: y = 16'b0000101101010000;
        3: y = 16'b0001000011101111;
        4: y = 16'b0001011010000100;
        5: y = 16'b0001110000001011;
        6: y = 16'b0010000110000000;
        7: y = 16'b0010011011100001;
        8: y = 16'b0010110000101010;
        9: y = 16'b0011000101011000;
        10: y = 16'b0011011001100111;
        11: y = 16'b0011101101010101;
        12: y = 16'b0100000000011110;
        13: y = 16'b0100010010111111;
        14: y = 16'b0100100100110111;
        15: y = 16'b0100110110000001;
        16: y = 16'b0101000110011011;
        17: y = 16'b0101010110000011;
        18: y = 16'b0101100100110110;
        19: y = 16'b0101110010110010;
        20: y = 16'b0101111111110101;
        21: y = 16'b0110001011111101;
        22: y = 16'b0110010111000111;
        23: y = 16'b0110100001010011;
        24: y = 16'b0110101010011111;
        25: y = 16'b0110110010101001;
        26: y = 16'b0110111001110000;
        27: y = 16'b0110111111110011;
        28: y = 16'b0111000100110000;
        29: y = 16'b0111001000101000;
        30: y = 16'b0111001011011010;
        31: y = 16'b0111001101000100;
        32: y = 16'b0111001101101000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=440.0Hz, Fs=52734Hz, 16-bit, Volume 15/15 bit

module table_52734_A
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 30;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000011000001010;
        2: y = 16'b0000110000010000;
        3: y = 16'b0001001000001110;
        4: y = 16'b0001011111111111;
        5: y = 16'b0001110111011111;
        6: y = 16'b0010001110101010;
        7: y = 16'b0010100101011100;
        8: y = 16'b0010111011110001;
        9: y = 16'b0011010001100101;
        10: y = 16'b0011100110110100;
        11: y = 16'b0011111011011011;
        12: y = 16'b0100001111010110;
        13: y = 16'b0100100010100001;
        14: y = 16'b0100110100111001;
        15: y = 16'b0101000110011011;
        16: y = 16'b0101010111000011;
        17: y = 16'b0101100110110000;
        18: y = 16'b0101110101011110;
        19: y = 16'b0110000011001010;
        20: y = 16'b0110001111110010;
        21: y = 16'b0110011011010100;
        22: y = 16'b0110100101101110;
        23: y = 16'b0110101110111110;
        24: y = 16'b0110110111000010;
        25: y = 16'b0110111101111001;
        26: y = 16'b0111000011100010;
        27: y = 16'b0111000111111100;
        28: y = 16'b0111001011000110;
        29: y = 16'b0111001101000000;
        30: y = 16'b0111001101101000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=466.16Hz, Fs=52734Hz, 16-bit, Volume 15/15 bit

module table_52734_As
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 28;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000011001111001;
        2: y = 16'b0000110011101100;
        3: y = 16'b0001001101010101;
        4: y = 16'b0001100110101110;
        5: y = 16'b0001111111110011;
        6: y = 16'b0010011000011110;
        7: y = 16'b0010110000101010;
        8: y = 16'b0011001000010011;
        9: y = 16'b0011011111010011;
        10: y = 16'b0011110101100110;
        11: y = 16'b0100001011001000;
        12: y = 16'b0100011111110100;
        13: y = 16'b0100110011100111;
        14: y = 16'b0101000110011011;
        15: y = 16'b0101011000001101;
        16: y = 16'b0101101000111010;
        17: y = 16'b0101111000011111;
        18: y = 16'b0110000110111000;
        19: y = 16'b0110010100000010;
        20: y = 16'b0110011111111010;
        21: y = 16'b0110101010011111;
        22: y = 16'b0110110011101110;
        23: y = 16'b0110111011100101;
        24: y = 16'b0111000010000011;
        25: y = 16'b0111000111000111;
        26: y = 16'b0111001010101110;
        27: y = 16'b0111001100111010;
        28: y = 16'b0111001101101000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=493.88Hz, Fs=52734Hz, 16-bit, Volume 15/15 bit

module table_52734_B
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 27;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000011010110110;
        2: y = 16'b0000110101100110;
        3: y = 16'b0001010000001010;
        4: y = 16'b0001101010011101;
        5: y = 16'b0010000100011001;
        6: y = 16'b0010011101111001;
        7: y = 16'b0010110110110110;
        8: y = 16'b0011001111001011;
        9: y = 16'b0011100110110100;
        10: y = 16'b0011111101101011;
        11: y = 16'b0100010011101010;
        12: y = 16'b0100101000101111;
        13: y = 16'b0100111100110010;
        14: y = 16'b0101001111110010;
        15: y = 16'b0101100001101000;
        16: y = 16'b0101110010010010;
        17: y = 16'b0110000001101100;
        18: y = 16'b0110001111110010;
        19: y = 16'b0110011100100001;
        20: y = 16'b0110100111111000;
        21: y = 16'b0110110001110010;
        22: y = 16'b0110111010001111;
        23: y = 16'b0111000001001100;
        24: y = 16'b0111000110100111;
        25: y = 16'b0111001010100000;
        26: y = 16'b0111001100110110;
        27: y = 16'b0111001101101000;
        default: y = 16'b0;
        endcase

endmodule

