`include "../arty_a7_35_pmod_mic3/board_specific_top.sv"
