`define FORCE_NO_INSTANTIATE_TM1638_BOARD_CONTROLLER_MODULE
`ifndef INSTANTIATE_GRAPHICS_INTERFACE_MODULE
`define VIRTUAL_TM1638_BOARD_CONTROLLER_GRAPHICS
`define INSTANTIATE_GRAPHICS_INTERFACE_MODULE
`endif
`include "../tang_nano_9k_hdmi_tm1638/board_specific_top.sv"
