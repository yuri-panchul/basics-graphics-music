//Copyright (C)2014-2025 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.11.03 Education
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9
//Device Version: C
//Created Time: Wed Dec 31 14:37:51 2025

module Gowin_pROM (dout, clk, oce, ce, reset, ad);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input [10:0] ad;

wire [23:0] prom_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[23:0],dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 8;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h0010387CFEFEFE6C7EFFE7C3FFDBFF7E7E8199BD81A5817E0000000000000000;
defparam prom_inst_0.INIT_RAM_01 = 256'h0000183C3C180000003810EEFE7C3810003C18E7FF183C3C0010387CFE7C3810;
defparam prom_inst_0.INIT_RAM_02 = 256'h78CCCCCC7D0F070FFFC399BDBD99C3FF003C664242663C00FFFFE7C3C3E7FFFF;
defparam prom_inst_0.INIT_RAM_03 = 256'h00105438EE3854101C0EE272161A141800F078080A0A0C08187E183C6666663C;
defparam prom_inst_0.INIT_RAM_04 = 256'h004400444444444400183C5A185A3C1800020E3EFE3E0E020080E0F8FEF8E080;
defparam prom_inst_0.INIT_RAM_05 = 256'h7E183C5A185A3C18007E7E0000000000708838444438221C001212121212927E;
defparam prom_inst_0.INIT_RAM_06 = 256'h00003060FE6030000000180CFE0C180000183C5A1818181800181818185A3C18;
defparam prom_inst_0.INIT_RAM_07 = 256'h000010387CFEFE000000FEFE7C38100000002442FF4224000000FEC0C0C00000;
defparam prom_inst_0.INIT_RAM_08 = 256'h004444FE44FE4444000000000000242400100010101010100000000000000000;
defparam prom_inst_0.INIT_RAM_09 = 256'h0000000000201010007A848A4830483000844A2450A844000010FC167CD07C10;
defparam prom_inst_0.INIT_RAM_0A = 256'h00002020F820200000006618FF18660000601008080810600018204040402018;
defparam prom_inst_0.INIT_RAM_0B = 256'h0080402010080402003000000000000000000000FC0000002010100000000000;
defparam prom_inst_0.INIT_RAM_0C = 256'h007C82023C02827C00FE80807C02827C007C101010503010007CC2A2928A867C;
defparam prom_inst_0.INIT_RAM_0D = 256'h00202020100804FC007C8282FC80827C007C820202FC80FE000404FE8444241C;
defparam prom_inst_0.INIT_RAM_0E = 256'h20101000000010000000100000001000007C82027E82827C007C8282827C827C;
defparam prom_inst_0.INIT_RAM_0F = 256'h0020002010088478002010080408102000007E00007E00000008102040201008;
defparam prom_inst_0.INIT_RAM_10 = 256'h007C82808080827C00FC8282FC8282FC00828282FE82827C007C809EA29E827C;
defparam prom_inst_0.INIT_RAM_11 = 256'h007C828E8080827C00808080F88080FE00FE8080F88080FE00F88482828284F8;
defparam prom_inst_0.INIT_RAM_12 = 256'h00828488F09088840078848404040404007C10101010107C00828282FE828282;
defparam prom_inst_0.INIT_RAM_13 = 256'h007C82828282827C0082868A92A2C2820082828292AAC68200FE808080808080;
defparam prom_inst_0.INIT_RAM_14 = 256'h007C82027C80827C00828282FC8282FC007C8A928282827C00808080FC8282FC;
defparam prom_inst_0.INIT_RAM_15 = 256'h0082C6AA928282820010284482828282007C82828282828200101010101010FE;
defparam prom_inst_0.INIT_RAM_16 = 256'h007840404040407800FE4020100804FE00101010284482820082442810284482;
defparam prom_inst_0.INIT_RAM_17 = 256'hFF00000000000000000000008244281000780808080808780002040810204080;
defparam prom_inst_0.INIT_RAM_18 = 256'h007C8280827C0000007C42427C404040007CC47C047800000000000000102030;
defparam prom_inst_0.INIT_RAM_19 = 256'h78047C84847C0000002020202038201C007C80F884780000007C84847C040404;
defparam prom_inst_0.INIT_RAM_1A = 256'h0044487048444040304808080808000800381010103000100044444478404040;
defparam prom_inst_0.INIT_RAM_1B = 256'h007C8282827C000000444444447800000092929292EC0000000C101010101010;
defparam prom_inst_0.INIT_RAM_1C = 256'h00FC027C807C0000004040404038000006047C84847C000040407C42427C0000;
defparam prom_inst_0.INIT_RAM_1D = 256'h006C929292820000001028444444000000788484848400000018202020702020;
defparam prom_inst_0.INIT_RAM_1E = 256'h000E10103010100E00FC402010FC0000F8047C84848400000044281028440000;
defparam prom_inst_0.INIT_RAM_1F = 256'h00FE8282442810000000000000009C7200E01010181010E00000101010101010;
defparam prom_inst_0.INIT_RAM_20 = 256'h0076CC7C0C38827C007CC0FEC67C100E0076CCCCCCCC00CC70187CC6C0C0C67C;
defparam prom_inst_0.INIT_RAM_21 = 256'h70187CC0C07C00000076CC7C0C7830300076CC7C0C7810E00076CC7C0C7800CC;
defparam prom_inst_0.INIT_RAM_22 = 256'h003C181818380066007CC0FEC67C10E0007CC0FEC67C00C6007CC0FEC67C827C;
defparam prom_inst_0.INIT_RAM_23 = 256'h00C6C6FEC67C383800C6C6FEC67C00C6003C1818183810E0003C18181838827C;
defparam prom_inst_0.INIT_RAM_24 = 256'h000000F0808080F0000000F090E090E00000009090F0906000FE607860FE100E;
defparam prom_inst_0.INIT_RAM_25 = 256'h0076CCCCCCCC10E00076CCCCCCCC827C007CC6C6C67C10E0007CC6C6C67C00C6;
defparam prom_inst_0.INIT_RAM_26 = 256'h00187CD6D0D67C18007CC6C6C6C600C6007CC6C6C6C67CC6F80C7CCCCCCC00CC;
defparam prom_inst_0.INIT_RAM_27 = 256'h70D818183C181B0E06CCDECCC4F8CCF800187E187E183C6600DCF260F0606C38;
defparam prom_inst_0.INIT_RAM_28 = 256'h0076CCCCCCCC100E007CC6C6C67C100E003C18181838100E0076CC7C0C78100E;
defparam prom_inst_0.INIT_RAM_29 = 256'h00007C00386C6C3800007E00343C0C3800C6CEDEF6E698660066666666DC9866;
defparam prom_inst_0.INIT_RAM_2A = 256'h001E8C46FED0C8C000000C0CFC0000000000C0C0FC000000007CC6C660300030;
defparam prom_inst_0.INIT_RAM_2B = 256'h0000D86C366CD8000000366CD86C360000183C3C18180018000CBE5CECD0C8C0;
defparam prom_inst_0.INIT_RAM_2C = 256'h000000E080E00000000000E0A0E08080000000E0A0E020E08822882288228822;
defparam prom_inst_0.INIT_RAM_2D = 256'h363636FE000000000000004040E04060000000E0C0A0C000000000E0A0E02020;
defparam prom_inst_0.INIT_RAM_2E = 256'h363636F606FE00003636363636363636363636F606F63636181818F818F80000;
defparam prom_inst_0.INIT_RAM_2F = 256'h181818F800000000000000F818F81818000000FE36363636000000FE06F63636;
defparam prom_inst_0.INIT_RAM_30 = 256'h1818181F18181818181818FF00000000000000FF181818180000001F18181818;
defparam prom_inst_0.INIT_RAM_31 = 256'h36363637363636361818181F181F1818181818FF18181818000000FF00000000;
defparam prom_inst_0.INIT_RAM_32 = 256'h363636F700FF0000000000FF00F7363636363637303F00000000003F30373636;
defparam prom_inst_0.INIT_RAM_33 = 256'h000000FF00FF1818363636F700F73636000000FF00FF00003636363730373636;
defparam prom_inst_0.INIT_RAM_34 = 256'h0000003F36363636363636FF00000000181818FF00FF0000000000FF36363636;
defparam prom_inst_0.INIT_RAM_35 = 256'h363636FF363636363636363F000000001818181F181F00000000001F181F1818;
defparam prom_inst_0.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFF1818181F00000000000000F818181818181818FF18FF1818;
defparam prom_inst_0.INIT_RAM_37 = 256'h00000000FFFFFFFF0F0F0F0F0F0F0F0FF0F0F0F0F0F0F0F0FFFFFFFF00000000;
defparam prom_inst_0.INIT_RAM_38 = 256'h00486C6CEC7E020000F06060606062FE40DCC6C6CCD8CC780076DCC8CC740000;
defparam prom_inst_0.INIT_RAM_39 = 256'h00101818D87E000080F8CCCCCCCC00000070C8C8D07E000000FE6230183062FE;
defparam prom_inst_0.INIT_RAM_3A = 256'h0078CCCC7C18223C00EE286CC6C6C67C007CC6C6FEC6C67C38107CD6D67C1038;
defparam prom_inst_0.INIT_RAM_3B = 256'h00C6C6C6C6C67C00007CC0F8C07C000000C07CF29E7C06000000669999660000;
defparam prom_inst_0.INIT_RAM_3C = 256'h007C001830603018007C0030180C1830007E0018187E18180000FE00FE00FE00;
defparam prom_inst_0.INIT_RAM_3D = 256'h0000DC7600DC7600000018007E00180070D8D8181818181818181818181B1B0E;
defparam prom_inst_0.INIT_RAM_3E = 256'h003C6CEC0C0C0C0F000000180000000000000018180000000000000000386C38;
defparam prom_inst_0.INIT_RAM_3F = 256'h000000000000000000003C3C3C3C000000000000F0C030F0000000006C6C6CD8;

endmodule //Gowin_pROM
