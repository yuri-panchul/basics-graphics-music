`define USE_DIGILENT_PMOD_MIC3
`include "../saylinx/board_specific_top.sv"
