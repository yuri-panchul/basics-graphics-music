`include "config.svh"

module lab_top
# (
    parameter  clk_mhz       = 50,
               w_key         = 4,
               w_sw          = 8,
               w_led         = 8,
               w_digit       = 8,
               w_gpio        = 100,

               screen_width  = 640,
               screen_height = 480,

               w_red         = 4,
               w_green       = 4,
               w_blue        = 4,

               w_x           = $clog2 ( screen_width  ),
               w_y           = $clog2 ( screen_height )
)
(
    input                        clk,
    input                        slow_clk,
    input                        rst,

    // Keys, switches, LEDs

    input        [w_key   - 1:0] key,
    input        [w_sw    - 1:0] sw,
    output logic [w_led   - 1:0] led,

    // A dynamic seven-segment display

    output logic [          7:0] abcdefgh,
    output logic [w_digit - 1:0] digit,

    // Graphics

    input        [w_x     - 1:0] x,
    input        [w_y     - 1:0] y,

    output logic [w_red   - 1:0] red,
    output logic [w_green - 1:0] green,
    output logic [w_blue  - 1:0] blue,

    // Microphone, sound output and UART

    input        [         23:0] mic,
    output       [         15:0] sound,

    input                        uart_rx,
    output                       uart_tx,

    // General-purpose Input/Output

    inout        [w_gpio  - 1:0] gpio
);

    //------------------------------------------------------------------------

       assign led        = '0;
       assign abcdefgh   = '0;
       assign digit      = '0;
    // assign red        = '0;
    // assign green      = '0;
    // assign blue       = '0;
       assign sound      = '0;
       assign uart_tx    = '1;

    //------------------------------------------------------------------------
    // Pattern 1

    /**/

    always_comb
    begin
        red   = '0;
        green = '0;
        blue  = '0;

        if(x < screen_width && y < screen_height)
        begin

            if (x < 128)
            begin
                red = x[w_red+3:3];
            end
    
            if (x >= 128 && x < 128+128)
            begin
                green = x[w_green+3:3];
            end
    
            if (x >= 128+128 && x < 128+128+128)
            begin
                blue = x[w_blue+3:3];
            end
    
            if (x >= 128+128+128 && x < 128+128+128+128)
            begin
                red = x[w_red+3:3];
                green = x[w_green+3:3];
            end
    
            if (x >= 128+128+128+128 && x < 128+128+128+128+128)
            begin
                green = x[6:3];
                blue = x[6:3];
            end

        end
    end
    
endmodule
