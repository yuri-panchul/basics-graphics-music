`define USE_DIGILENT_PMOD_MIC3
`include "../saylinx_pmod_mic3/board_specific_top.sv"
