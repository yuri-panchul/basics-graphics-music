// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=261.63Hz, Fs=48828Hz, 16-bit, Volume 14/15 bit

module table_48828_C
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 47;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001000100011;
        2: y = 16'b0000010001000110;
        3: y = 16'b0000011001101000;
        4: y = 16'b0000100010001000;
        5: y = 16'b0000101010100101;
        6: y = 16'b0000110010111111;
        7: y = 16'b0000111011010110;
        8: y = 16'b0001000011101000;
        9: y = 16'b0001001011110110;
        10: y = 16'b0001010011111110;
        11: y = 16'b0001011100000000;
        12: y = 16'b0001100011111011;
        13: y = 16'b0001101011110000;
        14: y = 16'b0001110011011100;
        15: y = 16'b0001111011000001;
        16: y = 16'b0010000010011101;
        17: y = 16'b0010001001101111;
        18: y = 16'b0010010000110111;
        19: y = 16'b0010010111110101;
        20: y = 16'b0010011110101001;
        21: y = 16'b0010100101010001;
        22: y = 16'b0010101011101101;
        23: y = 16'b0010110001111101;
        24: y = 16'b0010111000000000;
        25: y = 16'b0010111101110110;
        26: y = 16'b0011000011011110;
        27: y = 16'b0011001000111001;
        28: y = 16'b0011001110000101;
        29: y = 16'b0011010011000010;
        30: y = 16'b0011010111110000;
        31: y = 16'b0011011100001111;
        32: y = 16'b0011100000011110;
        33: y = 16'b0011100100011101;
        34: y = 16'b0011101000001100;
        35: y = 16'b0011101011101010;
        36: y = 16'b0011101110110111;
        37: y = 16'b0011110001110100;
        38: y = 16'b0011110100011110;
        39: y = 16'b0011110110111000;
        40: y = 16'b0011111001000000;
        41: y = 16'b0011111010110110;
        42: y = 16'b0011111100011010;
        43: y = 16'b0011111101101100;
        44: y = 16'b0011111110101100;
        45: y = 16'b0011111111011001;
        46: y = 16'b0011111111110101;
        47: y = 16'b0011111111111110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=277.18Hz, Fs=48828Hz, 16-bit, Volume 14/15 bit

module table_48828_Cs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 44;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001001001001;
        2: y = 16'b0000010010010001;
        3: y = 16'b0000011011010111;
        4: y = 16'b0000100100011011;
        5: y = 16'b0000101101011101;
        6: y = 16'b0000110110011010;
        7: y = 16'b0000111111010011;
        8: y = 16'b0001001000000111;
        9: y = 16'b0001010000110101;
        10: y = 16'b0001011001011101;
        11: y = 16'b0001100001111101;
        12: y = 16'b0001101010010101;
        13: y = 16'b0001110010100101;
        14: y = 16'b0001111010101011;
        15: y = 16'b0010000010100111;
        16: y = 16'b0010001010011001;
        17: y = 16'b0010010001111111;
        18: y = 16'b0010011001011001;
        19: y = 16'b0010100000100111;
        20: y = 16'b0010100111101000;
        21: y = 16'b0010101110011011;
        22: y = 16'b0010110101000000;
        23: y = 16'b0010111011010110;
        24: y = 16'b0011000001011101;
        25: y = 16'b0011000111010100;
        26: y = 16'b0011001100111010;
        27: y = 16'b0011010010010001;
        28: y = 16'b0011010111010101;
        29: y = 16'b0011011100001001;
        30: y = 16'b0011100000101010;
        31: y = 16'b0011100100111001;
        32: y = 16'b0011101000110110;
        33: y = 16'b0011101100011111;
        34: y = 16'b0011101111110101;
        35: y = 16'b0011110010111000;
        36: y = 16'b0011110101100110;
        37: y = 16'b0011111000000001;
        38: y = 16'b0011111010001000;
        39: y = 16'b0011111011111010;
        40: y = 16'b0011111101010111;
        41: y = 16'b0011111110100000;
        42: y = 16'b0011111111010100;
        43: y = 16'b0011111111110100;
        44: y = 16'b0011111111111110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=293.66Hz, Fs=48828Hz, 16-bit, Volume 14/15 bit

module table_48828_D
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 42;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001001100101;
        2: y = 16'b0000010011001000;
        3: y = 16'b0000011100101010;
        4: y = 16'b0000100110001010;
        5: y = 16'b0000101111100110;
        6: y = 16'b0000111000111101;
        7: y = 16'b0001000010010000;
        8: y = 16'b0001001011011101;
        9: y = 16'b0001010100100011;
        10: y = 16'b0001011101100001;
        11: y = 16'b0001100110010111;
        12: y = 16'b0001101111000100;
        13: y = 16'b0001110111100111;
        14: y = 16'b0001111111111111;
        15: y = 16'b0010001000001100;
        16: y = 16'b0010010000001100;
        17: y = 16'b0010011000000000;
        18: y = 16'b0010011111100110;
        19: y = 16'b0010100110111110;
        20: y = 16'b0010101110000111;
        21: y = 16'b0010110101000000;
        22: y = 16'b0010111011101001;
        23: y = 16'b0011000010000001;
        24: y = 16'b0011001000001000;
        25: y = 16'b0011001101111101;
        26: y = 16'b0011010011011111;
        27: y = 16'b0011011000101111;
        28: y = 16'b0011011101101011;
        29: y = 16'b0011100010010100;
        30: y = 16'b0011100110101000;
        31: y = 16'b0011101010100111;
        32: y = 16'b0011101110010010;
        33: y = 16'b0011110001100111;
        34: y = 16'b0011110100100110;
        35: y = 16'b0011110111010000;
        36: y = 16'b0011111001100011;
        37: y = 16'b0011111011100000;
        38: y = 16'b0011111101000111;
        39: y = 16'b0011111110010111;
        40: y = 16'b0011111111010000;
        41: y = 16'b0011111111110011;
        42: y = 16'b0011111111111110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=311.13Hz, Fs=48828Hz, 16-bit, Volume 14/15 bit

module table_48828_Ds
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 39;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001010010100;
        2: y = 16'b0000010100100110;
        3: y = 16'b0000011110110111;
        4: y = 16'b0000101001000100;
        5: y = 16'b0000110011001101;
        6: y = 16'b0000111101010000;
        7: y = 16'b0001000111001110;
        8: y = 16'b0001010001000100;
        9: y = 16'b0001011010110001;
        10: y = 16'b0001100100010101;
        11: y = 16'b0001101101101111;
        12: y = 16'b0001110110111101;
        13: y = 16'b0001111111111111;
        14: y = 16'b0010001000110100;
        15: y = 16'b0010010001011010;
        16: y = 16'b0010011001110001;
        17: y = 16'b0010100001111001;
        18: y = 16'b0010101001101111;
        19: y = 16'b0010110001010100;
        20: y = 16'b0010111000100111;
        21: y = 16'b0010111111100110;
        22: y = 16'b0011000110010010;
        23: y = 16'b0011001100101000;
        24: y = 16'b0011010010101010;
        25: y = 16'b0011011000010110;
        26: y = 16'b0011011101101011;
        27: y = 16'b0011100010101010;
        28: y = 16'b0011100111010000;
        29: y = 16'b0011101011011111;
        30: y = 16'b0011101111010101;
        31: y = 16'b0011110010110011;
        32: y = 16'b0011110101110111;
        33: y = 16'b0011111000100010;
        34: y = 16'b0011111010110011;
        35: y = 16'b0011111100101010;
        36: y = 16'b0011111110000111;
        37: y = 16'b0011111111001001;
        38: y = 16'b0011111111110001;
        39: y = 16'b0011111111111110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=329.63Hz, Fs=48828Hz, 16-bit, Volume 14/15 bit

module table_48828_E
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 37;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001010110111;
        2: y = 16'b0000010101101101;
        3: y = 16'b0000100000100001;
        4: y = 16'b0000101011010001;
        5: y = 16'b0000110101111011;
        6: y = 16'b0001000000100000;
        7: y = 16'b0001001010111101;
        8: y = 16'b0001010101010001;
        9: y = 16'b0001011111011100;
        10: y = 16'b0001101001011100;
        11: y = 16'b0001110011001111;
        12: y = 16'b0001111100110101;
        13: y = 16'b0010000110001101;
        14: y = 16'b0010001111010110;
        15: y = 16'b0010011000001101;
        16: y = 16'b0010100000110011;
        17: y = 16'b0010101001000111;
        18: y = 16'b0010110001000111;
        19: y = 16'b0010111000110011;
        20: y = 16'b0011000000001010;
        21: y = 16'b0011000111001010;
        22: y = 16'b0011001101110011;
        23: y = 16'b0011010100000101;
        24: y = 16'b0011011001111110;
        25: y = 16'b0011011111011110;
        26: y = 16'b0011100100100100;
        27: y = 16'b0011101001010000;
        28: y = 16'b0011101101100001;
        29: y = 16'b0011110001010110;
        30: y = 16'b0011110100110000;
        31: y = 16'b0011110111101101;
        32: y = 16'b0011111010001110;
        33: y = 16'b0011111100010010;
        34: y = 16'b0011111101111001;
        35: y = 16'b0011111111000011;
        36: y = 16'b0011111111101111;
        37: y = 16'b0011111111111110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=349.23Hz, Fs=48828Hz, 16-bit, Volume 14/15 bit

module table_48828_F
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 35;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001011011111;
        2: y = 16'b0000010110111100;
        3: y = 16'b0000100010010111;
        4: y = 16'b0000101101101101;
        5: y = 16'b0000111000111101;
        6: y = 16'b0001000100000110;
        7: y = 16'b0001001111000110;
        8: y = 16'b0001011001111100;
        9: y = 16'b0001100100100111;
        10: y = 16'b0001101111000100;
        11: y = 16'b0001111001010011;
        12: y = 16'b0010000011010010;
        13: y = 16'b0010001101000001;
        14: y = 16'b0010010110011101;
        15: y = 16'b0010011111100110;
        16: y = 16'b0010101000011010;
        17: y = 16'b0010110000111001;
        18: y = 16'b0010111001000001;
        19: y = 16'b0011000000110001;
        20: y = 16'b0011001000001000;
        21: y = 16'b0011001111000101;
        22: y = 16'b0011010101101000;
        23: y = 16'b0011011011101111;
        24: y = 16'b0011100001011010;
        25: y = 16'b0011100110101000;
        26: y = 16'b0011101011011000;
        27: y = 16'b0011101111101001;
        28: y = 16'b0011110011011100;
        29: y = 16'b0011110110110000;
        30: y = 16'b0011111001100011;
        31: y = 16'b0011111011110111;
        32: y = 16'b0011111101101010;
        33: y = 16'b0011111110111100;
        34: y = 16'b0011111111101110;
        35: y = 16'b0011111111111110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=369.99Hz, Fs=48828Hz, 16-bit, Volume 14/15 bit

module table_48828_Fs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 33;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001100001011;
        2: y = 16'b0000011000010101;
        3: y = 16'b0000100100011011;
        4: y = 16'b0000110000011100;
        5: y = 16'b0000111100010110;
        6: y = 16'b0001001000000111;
        7: y = 16'b0001010011101110;
        8: y = 16'b0001011111001001;
        9: y = 16'b0001101010010101;
        10: y = 16'b0001110101010011;
        11: y = 16'b0001111111111111;
        12: y = 16'b0010001010011001;
        13: y = 16'b0010010100011110;
        14: y = 16'b0010011110001111;
        15: y = 16'b0010100111101000;
        16: y = 16'b0010110000101001;
        17: y = 16'b0010111001010000;
        18: y = 16'b0011000001011101;
        19: y = 16'b0011001001001101;
        20: y = 16'b0011010000100000;
        21: y = 16'b0011010111010101;
        22: y = 16'b0011011101101011;
        23: y = 16'b0011100011100001;
        24: y = 16'b0011101000110110;
        25: y = 16'b0011101101101001;
        26: y = 16'b0011110001111001;
        27: y = 16'b0011110101100110;
        28: y = 16'b0011111000110000;
        29: y = 16'b0011111011010110;
        30: y = 16'b0011111101010111;
        31: y = 16'b0011111110110100;
        32: y = 16'b0011111111101011;
        33: y = 16'b0011111111111110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=392.0Hz, Fs=48828Hz, 16-bit, Volume 14/15 bit

module table_48828_G
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 31;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001100111110;
        2: y = 16'b0000011001111001;
        3: y = 16'b0000100110110001;
        4: y = 16'b0000110011100010;
        5: y = 16'b0001000000001010;
        6: y = 16'b0001001100101000;
        7: y = 16'b0001011000111010;
        8: y = 16'b0001100100111100;
        9: y = 16'b0001110000101111;
        10: y = 16'b0001111100001110;
        11: y = 16'b0010000111011001;
        12: y = 16'b0010010010001111;
        13: y = 16'b0010011100101100;
        14: y = 16'b0010100110101111;
        15: y = 16'b0010110000010111;
        16: y = 16'b0010111001100010;
        17: y = 16'b0011000010001110;
        18: y = 16'b0011001010011010;
        19: y = 16'b0011010010000110;
        20: y = 16'b0011011001001110;
        21: y = 16'b0011011111110100;
        22: y = 16'b0011100101110100;
        23: y = 16'b0011101011001110;
        24: y = 16'b0011110000000010;
        25: y = 16'b0011110100001111;
        26: y = 16'b0011110111110011;
        27: y = 16'b0011111010101111;
        28: y = 16'b0011111101000001;
        29: y = 16'b0011111110101010;
        30: y = 16'b0011111111101001;
        31: y = 16'b0011111111111110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=415.3Hz, Fs=48828Hz, 16-bit, Volume 14/15 bit

module table_48828_Gs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 29;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001101110111;
        2: y = 16'b0000011011101011;
        3: y = 16'b0000101001011010;
        4: y = 16'b0000110111000010;
        5: y = 16'b0001000100011111;
        6: y = 16'b0001010001101111;
        7: y = 16'b0001011110110000;
        8: y = 16'b0001101011011111;
        9: y = 16'b0001110111111001;
        10: y = 16'b0010000011111110;
        11: y = 16'b0010001111101001;
        12: y = 16'b0010011010111010;
        13: y = 16'b0010100101101101;
        14: y = 16'b0010110000000010;
        15: y = 16'b0010111001110101;
        16: y = 16'b0011000011000110;
        17: y = 16'b0011001011110010;
        18: y = 16'b0011010011110111;
        19: y = 16'b0011011011010101;
        20: y = 16'b0011100010001010;
        21: y = 16'b0011101000010100;
        22: y = 16'b0011101101110010;
        23: y = 16'b0011110010100100;
        24: y = 16'b0011110110101001;
        25: y = 16'b0011111001111111;
        26: y = 16'b0011111100100110;
        27: y = 16'b0011111110011110;
        28: y = 16'b0011111111100110;
        29: y = 16'b0011111111111110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=440.0Hz, Fs=48828Hz, 16-bit, Volume 14/15 bit

module table_48828_A
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 28;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001110010111;
        2: y = 16'b0000011100101010;
        3: y = 16'b0000101010111000;
        4: y = 16'b0000111000111101;
        5: y = 16'b0001000110110111;
        6: y = 16'b0001010100100011;
        7: y = 16'b0001100001111101;
        8: y = 16'b0001101111000100;
        9: y = 16'b0001111011110100;
        10: y = 16'b0010001000001100;
        11: y = 16'b0010010100001000;
        12: y = 16'b0010011111100110;
        13: y = 16'b0010101010100100;
        14: y = 16'b0010110101000000;
        15: y = 16'b0010111110110111;
        16: y = 16'b0011001000001000;
        17: y = 16'b0011010000110001;
        18: y = 16'b0011011000101111;
        19: y = 16'b0011100000000010;
        20: y = 16'b0011100110101000;
        21: y = 16'b0011101100011111;
        22: y = 16'b0011110001100111;
        23: y = 16'b0011110101111110;
        24: y = 16'b0011111001100011;
        25: y = 16'b0011111100010111;
        26: y = 16'b0011111110010111;
        27: y = 16'b0011111111100100;
        28: y = 16'b0011111111111110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=466.16Hz, Fs=48828Hz, 16-bit, Volume 14/15 bit

module table_48828_As
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 26;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001111011101;
        2: y = 16'b0000011110110111;
        3: y = 16'b0000101110001001;
        4: y = 16'b0000111101010000;
        5: y = 16'b0001001100001010;
        6: y = 16'b0001011010110001;
        7: y = 16'b0001101001000011;
        8: y = 16'b0001110110111101;
        9: y = 16'b0010000100011011;
        10: y = 16'b0010010001011010;
        11: y = 16'b0010011101110111;
        12: y = 16'b0010101001101111;
        13: y = 16'b0010110101000000;
        14: y = 16'b0010111111100110;
        15: y = 16'b0011001001100000;
        16: y = 16'b0011010010101010;
        17: y = 16'b0011011011000011;
        18: y = 16'b0011100010101010;
        19: y = 16'b0011101001011011;
        20: y = 16'b0011101111010101;
        21: y = 16'b0011110100011000;
        22: y = 16'b0011111000100010;
        23: y = 16'b0011111011110010;
        24: y = 16'b0011111110000111;
        25: y = 16'b0011111111100000;
        26: y = 16'b0011111111111110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=493.88Hz, Fs=48828Hz, 16-bit, Volume 14/15 bit

module table_48828_B
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 25;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000010000000101;
        2: y = 16'b0000100000000101;
        3: y = 16'b0000101111111110;
        4: y = 16'b0000111111101010;
        5: y = 16'b0001001111000110;
        6: y = 16'b0001011110001111;
        7: y = 16'b0001101100111111;
        8: y = 16'b0001111011010100;
        9: y = 16'b0010001001001010;
        10: y = 16'b0010010110011101;
        11: y = 16'b0010100011001010;
        12: y = 16'b0010101111001110;
        13: y = 16'b0010111010100110;
        14: y = 16'b0011000101001111;
        15: y = 16'b0011001111000101;
        16: y = 16'b0011011000001000;
        17: y = 16'b0011100000010100;
        18: y = 16'b0011100111100111;
        19: y = 16'b0011101110000000;
        20: y = 16'b0011110011011100;
        21: y = 16'b0011110111111011;
        22: y = 16'b0011111011011100;
        23: y = 16'b0011111101111101;
        24: y = 16'b0011111111011110;
        25: y = 16'b0011111111111110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=261.63Hz, Fs=64453Hz, 16-bit, Volume 14/15 bit

module table_64453_C
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 62;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000000110011111;
        2: y = 16'b0000001100111110;
        3: y = 16'b0000010011011100;
        4: y = 16'b0000011001111001;
        5: y = 16'b0000100000010110;
        6: y = 16'b0000100110110001;
        7: y = 16'b0000101101001010;
        8: y = 16'b0000110011100010;
        9: y = 16'b0000111001110111;
        10: y = 16'b0001000000001010;
        11: y = 16'b0001000110011011;
        12: y = 16'b0001001100101000;
        13: y = 16'b0001010010110011;
        14: y = 16'b0001011000111010;
        15: y = 16'b0001011110111101;
        16: y = 16'b0001100100111100;
        17: y = 16'b0001101010111000;
        18: y = 16'b0001110000101111;
        19: y = 16'b0001110110100001;
        20: y = 16'b0001111100001110;
        21: y = 16'b0010000001110111;
        22: y = 16'b0010000111011001;
        23: y = 16'b0010001100110111;
        24: y = 16'b0010010010001111;
        25: y = 16'b0010010111100000;
        26: y = 16'b0010011100101100;
        27: y = 16'b0010100001110000;
        28: y = 16'b0010100110101111;
        29: y = 16'b0010101011100110;
        30: y = 16'b0010110000010111;
        31: y = 16'b0010110101000000;
        32: y = 16'b0010111001100010;
        33: y = 16'b0010111101111100;
        34: y = 16'b0011000010001110;
        35: y = 16'b0011000110011000;
        36: y = 16'b0011001010011010;
        37: y = 16'b0011001110010100;
        38: y = 16'b0011010010000110;
        39: y = 16'b0011010101101111;
        40: y = 16'b0011011001001110;
        41: y = 16'b0011011100100110;
        42: y = 16'b0011011111110100;
        43: y = 16'b0011100010111000;
        44: y = 16'b0011100101110100;
        45: y = 16'b0011101000100110;
        46: y = 16'b0011101011001110;
        47: y = 16'b0011101101101101;
        48: y = 16'b0011110000000010;
        49: y = 16'b0011110010001101;
        50: y = 16'b0011110100001111;
        51: y = 16'b0011110110000110;
        52: y = 16'b0011110111110011;
        53: y = 16'b0011111001010110;
        54: y = 16'b0011111010101111;
        55: y = 16'b0011111011111101;
        56: y = 16'b0011111101000001;
        57: y = 16'b0011111101111011;
        58: y = 16'b0011111110101010;
        59: y = 16'b0011111111001111;
        60: y = 16'b0011111111101001;
        61: y = 16'b0011111111111001;
        62: y = 16'b0011111111111110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=277.18Hz, Fs=64453Hz, 16-bit, Volume 14/15 bit

module table_64453_Cs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 58;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000000110111100;
        2: y = 16'b0000001101110111;
        3: y = 16'b0000010100110010;
        4: y = 16'b0000011011101011;
        5: y = 16'b0000100010100100;
        6: y = 16'b0000101001011010;
        7: y = 16'b0000110000001111;
        8: y = 16'b0000110111000010;
        9: y = 16'b0000111101110010;
        10: y = 16'b0001000100011111;
        11: y = 16'b0001001011001000;
        12: y = 16'b0001010001101111;
        13: y = 16'b0001011000010001;
        14: y = 16'b0001011110110000;
        15: y = 16'b0001100101001001;
        16: y = 16'b0001101011011111;
        17: y = 16'b0001110001101111;
        18: y = 16'b0001110111111001;
        19: y = 16'b0001111101111111;
        20: y = 16'b0010000011111110;
        21: y = 16'b0010001001110111;
        22: y = 16'b0010001111101001;
        23: y = 16'b0010010101010101;
        24: y = 16'b0010011010111010;
        25: y = 16'b0010100000010111;
        26: y = 16'b0010100101101101;
        27: y = 16'b0010101010111100;
        28: y = 16'b0010110000000010;
        29: y = 16'b0010110101000000;
        30: y = 16'b0010111001110101;
        31: y = 16'b0010111110100010;
        32: y = 16'b0011000011000110;
        33: y = 16'b0011000111100000;
        34: y = 16'b0011001011110010;
        35: y = 16'b0011001111111001;
        36: y = 16'b0011010011110111;
        37: y = 16'b0011010111101011;
        38: y = 16'b0011011011010101;
        39: y = 16'b0011011110110101;
        40: y = 16'b0011100010001010;
        41: y = 16'b0011100101010100;
        42: y = 16'b0011101000010100;
        43: y = 16'b0011101011001001;
        44: y = 16'b0011101101110010;
        45: y = 16'b0011110000010001;
        46: y = 16'b0011110010100100;
        47: y = 16'b0011110100101100;
        48: y = 16'b0011110110101001;
        49: y = 16'b0011111000011010;
        50: y = 16'b0011111001111111;
        51: y = 16'b0011111011011000;
        52: y = 16'b0011111100100110;
        53: y = 16'b0011111101101000;
        54: y = 16'b0011111110011110;
        55: y = 16'b0011111111001000;
        56: y = 16'b0011111111100110;
        57: y = 16'b0011111111111000;
        58: y = 16'b0011111111111110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=293.66Hz, Fs=64453Hz, 16-bit, Volume 14/15 bit

module table_64453_D
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 55;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000000111010100;
        2: y = 16'b0000001110100111;
        3: y = 16'b0000010101111010;
        4: y = 16'b0000011101001011;
        5: y = 16'b0000100100011011;
        6: y = 16'b0000101011101001;
        7: y = 16'b0000110010110101;
        8: y = 16'b0000111001111110;
        9: y = 16'b0001000001000101;
        10: y = 16'b0001001000000111;
        11: y = 16'b0001001111000110;
        12: y = 16'b0001010110000001;
        13: y = 16'b0001011100111000;
        14: y = 16'b0001100011101001;
        15: y = 16'b0001101010010101;
        16: y = 16'b0001110000111100;
        17: y = 16'b0001110111011101;
        18: y = 16'b0001111101111000;
        19: y = 16'b0010000100001100;
        20: y = 16'b0010001010011001;
        21: y = 16'b0010010000011111;
        22: y = 16'b0010010110011101;
        23: y = 16'b0010011100010100;
        24: y = 16'b0010100010000010;
        25: y = 16'b0010100111101000;
        26: y = 16'b0010101101000101;
        27: y = 16'b0010110010011001;
        28: y = 16'b0010110111100100;
        29: y = 16'b0010111100100101;
        30: y = 16'b0011000001011101;
        31: y = 16'b0011000110001010;
        32: y = 16'b0011001010101101;
        33: y = 16'b0011001111000101;
        34: y = 16'b0011010011010011;
        35: y = 16'b0011010111010101;
        36: y = 16'b0011011011001101;
        37: y = 16'b0011011110111001;
        38: y = 16'b0011100010011001;
        39: y = 16'b0011100101101101;
        40: y = 16'b0011101000110110;
        41: y = 16'b0011101011110010;
        42: y = 16'b0011101110100010;
        43: y = 16'b0011110001000101;
        44: y = 16'b0011110011011100;
        45: y = 16'b0011110101100110;
        46: y = 16'b0011110111100100;
        47: y = 16'b0011111001010100;
        48: y = 16'b0011111010111000;
        49: y = 16'b0011111100001110;
        50: y = 16'b0011111101010111;
        51: y = 16'b0011111110010011;
        52: y = 16'b0011111111000010;
        53: y = 16'b0011111111100011;
        54: y = 16'b0011111111110111;
        55: y = 16'b0011111111111110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=311.13Hz, Fs=64453Hz, 16-bit, Volume 14/15 bit

module table_64453_Ds
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 52;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000000111101111;
        2: y = 16'b0000001111011101;
        3: y = 16'b0000010111001011;
        4: y = 16'b0000011110110111;
        5: y = 16'b0000100110100001;
        6: y = 16'b0000101110001001;
        7: y = 16'b0000110101101110;
        8: y = 16'b0000111101010000;
        9: y = 16'b0001000100101111;
        10: y = 16'b0001001100001010;
        11: y = 16'b0001010011100000;
        12: y = 16'b0001011010110001;
        13: y = 16'b0001100001111101;
        14: y = 16'b0001101001000011;
        15: y = 16'b0001110000000100;
        16: y = 16'b0001110110111101;
        17: y = 16'b0001111101110000;
        18: y = 16'b0010000100011011;
        19: y = 16'b0010001010111111;
        20: y = 16'b0010010001011010;
        21: y = 16'b0010010111101101;
        22: y = 16'b0010011101110111;
        23: y = 16'b0010100011111000;
        24: y = 16'b0010101001101111;
        25: y = 16'b0010101111011101;
        26: y = 16'b0010110101000000;
        27: y = 16'b0010111010011000;
        28: y = 16'b0010111111100110;
        29: y = 16'b0011000100101001;
        30: y = 16'b0011001001100000;
        31: y = 16'b0011001110001011;
        32: y = 16'b0011010010101010;
        33: y = 16'b0011010110111101;
        34: y = 16'b0011011011000011;
        35: y = 16'b0011011110111101;
        36: y = 16'b0011100010101010;
        37: y = 16'b0011100110001001;
        38: y = 16'b0011101001011011;
        39: y = 16'b0011101100011111;
        40: y = 16'b0011101111010101;
        41: y = 16'b0011110001111110;
        42: y = 16'b0011110100011000;
        43: y = 16'b0011110110100100;
        44: y = 16'b0011111000100010;
        45: y = 16'b0011111010010001;
        46: y = 16'b0011111011110010;
        47: y = 16'b0011111101000011;
        48: y = 16'b0011111110000111;
        49: y = 16'b0011111110111011;
        50: y = 16'b0011111111100000;
        51: y = 16'b0011111111110111;
        52: y = 16'b0011111111111110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=329.63Hz, Fs=64453Hz, 16-bit, Volume 14/15 bit

module table_64453_E
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 49;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001000001101;
        2: y = 16'b0000010000011010;
        3: y = 16'b0000011000100101;
        4: y = 16'b0000100000101111;
        5: y = 16'b0000101000110111;
        6: y = 16'b0000110000111100;
        7: y = 16'b0000111000111101;
        8: y = 16'b0001000000111011;
        9: y = 16'b0001001000110101;
        10: y = 16'b0001010000101010;
        11: y = 16'b0001011000011010;
        12: y = 16'b0001100000000100;
        13: y = 16'b0001100111100111;
        14: y = 16'b0001101111000100;
        15: y = 16'b0001110110011001;
        16: y = 16'b0001111101100111;
        17: y = 16'b0010000100101100;
        18: y = 16'b0010001011101001;
        19: y = 16'b0010010010011100;
        20: y = 16'b0010011001000110;
        21: y = 16'b0010011111100110;
        22: y = 16'b0010100101111011;
        23: y = 16'b0010101100000110;
        24: y = 16'b0010110010000101;
        25: y = 16'b0010110111111000;
        26: y = 16'b0010111101011111;
        27: y = 16'b0011000010111010;
        28: y = 16'b0011001000001000;
        29: y = 16'b0011001101001001;
        30: y = 16'b0011010001111100;
        31: y = 16'b0011010110100010;
        32: y = 16'b0011011010111001;
        33: y = 16'b0011011111000010;
        34: y = 16'b0011100010111100;
        35: y = 16'b0011100110101000;
        36: y = 16'b0011101010000100;
        37: y = 16'b0011101101010001;
        38: y = 16'b0011110000001110;
        39: y = 16'b0011110010111011;
        40: y = 16'b0011110101011001;
        41: y = 16'b0011110111100110;
        42: y = 16'b0011111001100011;
        43: y = 16'b0011111011010000;
        44: y = 16'b0011111100101100;
        45: y = 16'b0011111101111000;
        46: y = 16'b0011111110110010;
        47: y = 16'b0011111111011100;
        48: y = 16'b0011111111110110;
        49: y = 16'b0011111111111110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=349.23Hz, Fs=64453Hz, 16-bit, Volume 14/15 bit

module table_64453_F
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 46;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001000101111;
        2: y = 16'b0000010001011110;
        3: y = 16'b0000011010001011;
        4: y = 16'b0000100010110111;
        5: y = 16'b0000101011011111;
        6: y = 16'b0000110100000101;
        7: y = 16'b0000111100100111;
        8: y = 16'b0001000101000100;
        9: y = 16'b0001001101011100;
        10: y = 16'b0001010101101110;
        11: y = 16'b0001011101111010;
        12: y = 16'b0001100101111111;
        13: y = 16'b0001101101111100;
        14: y = 16'b0001110101110001;
        15: y = 16'b0001111101011101;
        16: y = 16'b0010000101000000;
        17: y = 16'b0010001100011001;
        18: y = 16'b0010010011100111;
        19: y = 16'b0010011010101011;
        20: y = 16'b0010100001100010;
        21: y = 16'b0010101000001110;
        22: y = 16'b0010101110101110;
        23: y = 16'b0010110101000000;
        24: y = 16'b0010111011000101;
        25: y = 16'b0011000000111011;
        26: y = 16'b0011000110100100;
        27: y = 16'b0011001011111101;
        28: y = 16'b0011010001001000;
        29: y = 16'b0011010110000010;
        30: y = 16'b0011011010101101;
        31: y = 16'b0011011111001000;
        32: y = 16'b0011100011010001;
        33: y = 16'b0011100111001010;
        34: y = 16'b0011101010110010;
        35: y = 16'b0011101110001000;
        36: y = 16'b0011110001001100;
        37: y = 16'b0011110011111110;
        38: y = 16'b0011110110011111;
        39: y = 16'b0011111000101100;
        40: y = 16'b0011111010100111;
        41: y = 16'b0011111100010000;
        42: y = 16'b0011111101100101;
        43: y = 16'b0011111110101000;
        44: y = 16'b0011111111011000;
        45: y = 16'b0011111111110100;
        46: y = 16'b0011111111111110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=369.99Hz, Fs=64453Hz, 16-bit, Volume 14/15 bit

module table_64453_Fs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 44;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001001001001;
        2: y = 16'b0000010010010001;
        3: y = 16'b0000011011010111;
        4: y = 16'b0000100100011011;
        5: y = 16'b0000101101011101;
        6: y = 16'b0000110110011010;
        7: y = 16'b0000111111010011;
        8: y = 16'b0001001000000111;
        9: y = 16'b0001010000110101;
        10: y = 16'b0001011001011101;
        11: y = 16'b0001100001111101;
        12: y = 16'b0001101010010101;
        13: y = 16'b0001110010100101;
        14: y = 16'b0001111010101011;
        15: y = 16'b0010000010100111;
        16: y = 16'b0010001010011001;
        17: y = 16'b0010010001111111;
        18: y = 16'b0010011001011001;
        19: y = 16'b0010100000100111;
        20: y = 16'b0010100111101000;
        21: y = 16'b0010101110011011;
        22: y = 16'b0010110101000000;
        23: y = 16'b0010111011010110;
        24: y = 16'b0011000001011101;
        25: y = 16'b0011000111010100;
        26: y = 16'b0011001100111010;
        27: y = 16'b0011010010010001;
        28: y = 16'b0011010111010101;
        29: y = 16'b0011011100001001;
        30: y = 16'b0011100000101010;
        31: y = 16'b0011100100111001;
        32: y = 16'b0011101000110110;
        33: y = 16'b0011101100011111;
        34: y = 16'b0011101111110101;
        35: y = 16'b0011110010111000;
        36: y = 16'b0011110101100110;
        37: y = 16'b0011111000000001;
        38: y = 16'b0011111010001000;
        39: y = 16'b0011111011111010;
        40: y = 16'b0011111101010111;
        41: y = 16'b0011111110100000;
        42: y = 16'b0011111111010100;
        43: y = 16'b0011111111110100;
        44: y = 16'b0011111111111110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=392.0Hz, Fs=64453Hz, 16-bit, Volume 14/15 bit

module table_64453_G
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 41;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001001110011;
        2: y = 16'b0000010011100110;
        3: y = 16'b0000011101010111;
        4: y = 16'b0000100111000101;
        5: y = 16'b0000110000101111;
        6: y = 16'b0000111010010101;
        7: y = 16'b0001000011110101;
        8: y = 16'b0001001101001111;
        9: y = 16'b0001010110100001;
        10: y = 16'b0001011111101100;
        11: y = 16'b0001101000101101;
        12: y = 16'b0001110001100101;
        13: y = 16'b0001111010010010;
        14: y = 16'b0010000010110100;
        15: y = 16'b0010001011001001;
        16: y = 16'b0010010011010001;
        17: y = 16'b0010011011001011;
        18: y = 16'b0010100010110111;
        19: y = 16'b0010101010010011;
        20: y = 16'b0010110001100000;
        21: y = 16'b0010111000011100;
        22: y = 16'b0010111111000110;
        23: y = 16'b0011000101011111;
        24: y = 16'b0011001011100100;
        25: y = 16'b0011010001010111;
        26: y = 16'b0011010110110110;
        27: y = 16'b0011011100000001;
        28: y = 16'b0011100000111000;
        29: y = 16'b0011100101011001;
        30: y = 16'b0011101001100101;
        31: y = 16'b0011101101011010;
        32: y = 16'b0011110000111010;
        33: y = 16'b0011110100000011;
        34: y = 16'b0011110110110100;
        35: y = 16'b0011111001001111;
        36: y = 16'b0011111011010010;
        37: y = 16'b0011111100111110;
        38: y = 16'b0011111110010010;
        39: y = 16'b0011111111001110;
        40: y = 16'b0011111111110010;
        41: y = 16'b0011111111111110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=415.3Hz, Fs=64453Hz, 16-bit, Volume 14/15 bit

module table_64453_Gs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 39;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001010010100;
        2: y = 16'b0000010100100110;
        3: y = 16'b0000011110110111;
        4: y = 16'b0000101001000100;
        5: y = 16'b0000110011001101;
        6: y = 16'b0000111101010000;
        7: y = 16'b0001000111001110;
        8: y = 16'b0001010001000100;
        9: y = 16'b0001011010110001;
        10: y = 16'b0001100100010101;
        11: y = 16'b0001101101101111;
        12: y = 16'b0001110110111101;
        13: y = 16'b0001111111111111;
        14: y = 16'b0010001000110100;
        15: y = 16'b0010010001011010;
        16: y = 16'b0010011001110001;
        17: y = 16'b0010100001111001;
        18: y = 16'b0010101001101111;
        19: y = 16'b0010110001010100;
        20: y = 16'b0010111000100111;
        21: y = 16'b0010111111100110;
        22: y = 16'b0011000110010010;
        23: y = 16'b0011001100101000;
        24: y = 16'b0011010010101010;
        25: y = 16'b0011011000010110;
        26: y = 16'b0011011101101011;
        27: y = 16'b0011100010101010;
        28: y = 16'b0011100111010000;
        29: y = 16'b0011101011011111;
        30: y = 16'b0011101111010101;
        31: y = 16'b0011110010110011;
        32: y = 16'b0011110101110111;
        33: y = 16'b0011111000100010;
        34: y = 16'b0011111010110011;
        35: y = 16'b0011111100101010;
        36: y = 16'b0011111110000111;
        37: y = 16'b0011111111001001;
        38: y = 16'b0011111111110001;
        39: y = 16'b0011111111111110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=440.0Hz, Fs=64453Hz, 16-bit, Volume 14/15 bit

module table_64453_A
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 37;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001010110111;
        2: y = 16'b0000010101101101;
        3: y = 16'b0000100000100001;
        4: y = 16'b0000101011010001;
        5: y = 16'b0000110101111011;
        6: y = 16'b0001000000100000;
        7: y = 16'b0001001010111101;
        8: y = 16'b0001010101010001;
        9: y = 16'b0001011111011100;
        10: y = 16'b0001101001011100;
        11: y = 16'b0001110011001111;
        12: y = 16'b0001111100110101;
        13: y = 16'b0010000110001101;
        14: y = 16'b0010001111010110;
        15: y = 16'b0010011000001101;
        16: y = 16'b0010100000110011;
        17: y = 16'b0010101001000111;
        18: y = 16'b0010110001000111;
        19: y = 16'b0010111000110011;
        20: y = 16'b0011000000001010;
        21: y = 16'b0011000111001010;
        22: y = 16'b0011001101110011;
        23: y = 16'b0011010100000101;
        24: y = 16'b0011011001111110;
        25: y = 16'b0011011111011110;
        26: y = 16'b0011100100100100;
        27: y = 16'b0011101001010000;
        28: y = 16'b0011101101100001;
        29: y = 16'b0011110001010110;
        30: y = 16'b0011110100110000;
        31: y = 16'b0011110111101101;
        32: y = 16'b0011111010001110;
        33: y = 16'b0011111100010010;
        34: y = 16'b0011111101111001;
        35: y = 16'b0011111111000011;
        36: y = 16'b0011111111101111;
        37: y = 16'b0011111111111110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=466.16Hz, Fs=64453Hz, 16-bit, Volume 14/15 bit

module table_64453_As
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 35;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001011011111;
        2: y = 16'b0000010110111100;
        3: y = 16'b0000100010010111;
        4: y = 16'b0000101101101101;
        5: y = 16'b0000111000111101;
        6: y = 16'b0001000100000110;
        7: y = 16'b0001001111000110;
        8: y = 16'b0001011001111100;
        9: y = 16'b0001100100100111;
        10: y = 16'b0001101111000100;
        11: y = 16'b0001111001010011;
        12: y = 16'b0010000011010010;
        13: y = 16'b0010001101000001;
        14: y = 16'b0010010110011101;
        15: y = 16'b0010011111100110;
        16: y = 16'b0010101000011010;
        17: y = 16'b0010110000111001;
        18: y = 16'b0010111001000001;
        19: y = 16'b0011000000110001;
        20: y = 16'b0011001000001000;
        21: y = 16'b0011001111000101;
        22: y = 16'b0011010101101000;
        23: y = 16'b0011011011101111;
        24: y = 16'b0011100001011010;
        25: y = 16'b0011100110101000;
        26: y = 16'b0011101011011000;
        27: y = 16'b0011101111101001;
        28: y = 16'b0011110011011100;
        29: y = 16'b0011110110110000;
        30: y = 16'b0011111001100011;
        31: y = 16'b0011111011110111;
        32: y = 16'b0011111101101010;
        33: y = 16'b0011111110111100;
        34: y = 16'b0011111111101110;
        35: y = 16'b0011111111111110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=493.88Hz, Fs=64453Hz, 16-bit, Volume 14/15 bit

module table_64453_B
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 33;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001100001011;
        2: y = 16'b0000011000010101;
        3: y = 16'b0000100100011011;
        4: y = 16'b0000110000011100;
        5: y = 16'b0000111100010110;
        6: y = 16'b0001001000000111;
        7: y = 16'b0001010011101110;
        8: y = 16'b0001011111001001;
        9: y = 16'b0001101010010101;
        10: y = 16'b0001110101010011;
        11: y = 16'b0001111111111111;
        12: y = 16'b0010001010011001;
        13: y = 16'b0010010100011110;
        14: y = 16'b0010011110001111;
        15: y = 16'b0010100111101000;
        16: y = 16'b0010110000101001;
        17: y = 16'b0010111001010000;
        18: y = 16'b0011000001011101;
        19: y = 16'b0011001001001101;
        20: y = 16'b0011010000100000;
        21: y = 16'b0011010111010101;
        22: y = 16'b0011011101101011;
        23: y = 16'b0011100011100001;
        24: y = 16'b0011101000110110;
        25: y = 16'b0011101101101001;
        26: y = 16'b0011110001111001;
        27: y = 16'b0011110101100110;
        28: y = 16'b0011111000110000;
        29: y = 16'b0011111011010110;
        30: y = 16'b0011111101010111;
        31: y = 16'b0011111110110100;
        32: y = 16'b0011111111101011;
        33: y = 16'b0011111111111110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=261.63Hz, Fs=52734Hz, 16-bit, Volume 14/15 bit

module table_52734_C
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 50;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001000000011;
        2: y = 16'b0000010000000101;
        3: y = 16'b0000011000000110;
        4: y = 16'b0000100000000101;
        5: y = 16'b0000101000000011;
        6: y = 16'b0000101111111110;
        7: y = 16'b0000110111110110;
        8: y = 16'b0000111111101010;
        9: y = 16'b0001000111011010;
        10: y = 16'b0001001111000110;
        11: y = 16'b0001010110101101;
        12: y = 16'b0001011110001111;
        13: y = 16'b0001100101101010;
        14: y = 16'b0001101100111111;
        15: y = 16'b0001110100001101;
        16: y = 16'b0001111011010100;
        17: y = 16'b0010000010010011;
        18: y = 16'b0010001001001010;
        19: y = 16'b0010001111111000;
        20: y = 16'b0010010110011101;
        21: y = 16'b0010011100111001;
        22: y = 16'b0010100011001010;
        23: y = 16'b0010101001010010;
        24: y = 16'b0010101111001110;
        25: y = 16'b0010110101000000;
        26: y = 16'b0010111010100110;
        27: y = 16'b0011000000000000;
        28: y = 16'b0011000101001111;
        29: y = 16'b0011001010010000;
        30: y = 16'b0011001111000101;
        31: y = 16'b0011010011101101;
        32: y = 16'b0011011000001000;
        33: y = 16'b0011011100010101;
        34: y = 16'b0011100000010100;
        35: y = 16'b0011100100000100;
        36: y = 16'b0011100111100111;
        37: y = 16'b0011101010111011;
        38: y = 16'b0011101110000000;
        39: y = 16'b0011110000110110;
        40: y = 16'b0011110011011100;
        41: y = 16'b0011110101110100;
        42: y = 16'b0011110111111011;
        43: y = 16'b0011111001110011;
        44: y = 16'b0011111011011100;
        45: y = 16'b0011111100110100;
        46: y = 16'b0011111101111101;
        47: y = 16'b0011111110110101;
        48: y = 16'b0011111111011110;
        49: y = 16'b0011111111110110;
        50: y = 16'b0011111111111110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=277.18Hz, Fs=52734Hz, 16-bit, Volume 14/15 bit

module table_52734_Cs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 48;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001000011000;
        2: y = 16'b0000010000101111;
        3: y = 16'b0000011001000110;
        4: y = 16'b0000100001011010;
        5: y = 16'b0000101001101101;
        6: y = 16'b0000110001111100;
        7: y = 16'b0000111010001000;
        8: y = 16'b0001000010010000;
        9: y = 16'b0001001010010011;
        10: y = 16'b0001010010010010;
        11: y = 16'b0001011010001011;
        12: y = 16'b0001100001111101;
        13: y = 16'b0001101001101001;
        14: y = 16'b0001110001001110;
        15: y = 16'b0001111000101010;
        16: y = 16'b0001111111111111;
        17: y = 16'b0010000111001011;
        18: y = 16'b0010001110001101;
        19: y = 16'b0010010101000110;
        20: y = 16'b0010011011110101;
        21: y = 16'b0010100010011001;
        22: y = 16'b0010101000110001;
        23: y = 16'b0010101110111111;
        24: y = 16'b0010110101000000;
        25: y = 16'b0010111010110101;
        26: y = 16'b0011000000011101;
        27: y = 16'b0011000101110111;
        28: y = 16'b0011001011000101;
        29: y = 16'b0011010000000100;
        30: y = 16'b0011010100110101;
        31: y = 16'b0011011001011000;
        32: y = 16'b0011011101101011;
        33: y = 16'b0011100001110000;
        34: y = 16'b0011100101100101;
        35: y = 16'b0011101001001010;
        36: y = 16'b0011101100011111;
        37: y = 16'b0011101111100100;
        38: y = 16'b0011110010011001;
        39: y = 16'b0011110100111101;
        40: y = 16'b0011110111010000;
        41: y = 16'b0011111001010010;
        42: y = 16'b0011111011000011;
        43: y = 16'b0011111100100011;
        44: y = 16'b0011111101110010;
        45: y = 16'b0011111110101111;
        46: y = 16'b0011111111011011;
        47: y = 16'b0011111111110101;
        48: y = 16'b0011111111111110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=293.66Hz, Fs=52734Hz, 16-bit, Volume 14/15 bit

module table_52734_D
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 45;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001000111100;
        2: y = 16'b0000010001110111;
        3: y = 16'b0000011010110000;
        4: y = 16'b0000100011101000;
        5: y = 16'b0000101100011101;
        6: y = 16'b0000110101001110;
        7: y = 16'b0000111101111011;
        8: y = 16'b0001000110100011;
        9: y = 16'b0001001111000110;
        10: y = 16'b0001010111100011;
        11: y = 16'b0001011111111001;
        12: y = 16'b0001101000000111;
        13: y = 16'b0001110000001101;
        14: y = 16'b0001111000001011;
        15: y = 16'b0001111111111111;
        16: y = 16'b0010000111101001;
        17: y = 16'b0010001111001001;
        18: y = 16'b0010010110011101;
        19: y = 16'b0010011101100110;
        20: y = 16'b0010100100100010;
        21: y = 16'b0010101011010010;
        22: y = 16'b0010110001110100;
        23: y = 16'b0010111000001000;
        24: y = 16'b0010111110001110;
        25: y = 16'b0011000100000101;
        26: y = 16'b0011001001101101;
        27: y = 16'b0011001111000101;
        28: y = 16'b0011010100001101;
        29: y = 16'b0011011001000101;
        30: y = 16'b0011011101101011;
        31: y = 16'b0011100010000000;
        32: y = 16'b0011100110000100;
        33: y = 16'b0011101001110110;
        34: y = 16'b0011101101010101;
        35: y = 16'b0011110000100010;
        36: y = 16'b0011110011011100;
        37: y = 16'b0011110110000011;
        38: y = 16'b0011111000010111;
        39: y = 16'b0011111010011000;
        40: y = 16'b0011111100000101;
        41: y = 16'b0011111101011111;
        42: y = 16'b0011111110100100;
        43: y = 16'b0011111111010110;
        44: y = 16'b0011111111110100;
        45: y = 16'b0011111111111110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=311.13Hz, Fs=52734Hz, 16-bit, Volume 14/15 bit

module table_52734_Ds
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 42;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001001100101;
        2: y = 16'b0000010011001000;
        3: y = 16'b0000011100101010;
        4: y = 16'b0000100110001010;
        5: y = 16'b0000101111100110;
        6: y = 16'b0000111000111101;
        7: y = 16'b0001000010010000;
        8: y = 16'b0001001011011101;
        9: y = 16'b0001010100100011;
        10: y = 16'b0001011101100001;
        11: y = 16'b0001100110010111;
        12: y = 16'b0001101111000100;
        13: y = 16'b0001110111100111;
        14: y = 16'b0001111111111111;
        15: y = 16'b0010001000001100;
        16: y = 16'b0010010000001100;
        17: y = 16'b0010011000000000;
        18: y = 16'b0010011111100110;
        19: y = 16'b0010100110111110;
        20: y = 16'b0010101110000111;
        21: y = 16'b0010110101000000;
        22: y = 16'b0010111011101001;
        23: y = 16'b0011000010000001;
        24: y = 16'b0011001000001000;
        25: y = 16'b0011001101111101;
        26: y = 16'b0011010011011111;
        27: y = 16'b0011011000101111;
        28: y = 16'b0011011101101011;
        29: y = 16'b0011100010010100;
        30: y = 16'b0011100110101000;
        31: y = 16'b0011101010100111;
        32: y = 16'b0011101110010010;
        33: y = 16'b0011110001100111;
        34: y = 16'b0011110100100110;
        35: y = 16'b0011110111010000;
        36: y = 16'b0011111001100011;
        37: y = 16'b0011111011100000;
        38: y = 16'b0011111101000111;
        39: y = 16'b0011111110010111;
        40: y = 16'b0011111111010000;
        41: y = 16'b0011111111110011;
        42: y = 16'b0011111111111110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=329.63Hz, Fs=52734Hz, 16-bit, Volume 14/15 bit

module table_52734_E
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 40;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001010000011;
        2: y = 16'b0000010100000101;
        3: y = 16'b0000011110000101;
        4: y = 16'b0000101000000011;
        5: y = 16'b0000110001111100;
        6: y = 16'b0000111011110000;
        7: y = 16'b0001000101011111;
        8: y = 16'b0001001111000110;
        9: y = 16'b0001011000100110;
        10: y = 16'b0001100001111101;
        11: y = 16'b0001101011001010;
        12: y = 16'b0001110100001101;
        13: y = 16'b0001111101000101;
        14: y = 16'b0010000101110000;
        15: y = 16'b0010001110001101;
        16: y = 16'b0010010110011101;
        17: y = 16'b0010011110011110;
        18: y = 16'b0010100110001111;
        19: y = 16'b0010101101110000;
        20: y = 16'b0010110101000000;
        21: y = 16'b0010111011111110;
        22: y = 16'b0011000010101001;
        23: y = 16'b0011001001000001;
        24: y = 16'b0011001111000101;
        25: y = 16'b0011010100110101;
        26: y = 16'b0011011010010000;
        27: y = 16'b0011011111010101;
        28: y = 16'b0011100100000100;
        29: y = 16'b0011101000011101;
        30: y = 16'b0011101100011111;
        31: y = 16'b0011110000001001;
        32: y = 16'b0011110011011100;
        33: y = 16'b0011110110010111;
        34: y = 16'b0011111000111001;
        35: y = 16'b0011111011000011;
        36: y = 16'b0011111100110100;
        37: y = 16'b0011111110001100;
        38: y = 16'b0011111111001011;
        39: y = 16'b0011111111110001;
        40: y = 16'b0011111111111110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=349.23Hz, Fs=52734Hz, 16-bit, Volume 14/15 bit

module table_52734_F
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 38;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001010100101;
        2: y = 16'b0000010101001001;
        3: y = 16'b0000011111101010;
        4: y = 16'b0000101010001000;
        5: y = 16'b0000110100100010;
        6: y = 16'b0000111110110110;
        7: y = 16'b0001001001000010;
        8: y = 16'b0001010011000111;
        9: y = 16'b0001011101000011;
        10: y = 16'b0001100110110101;
        11: y = 16'b0001110000011011;
        12: y = 16'b0001111001110101;
        13: y = 16'b0010000011000010;
        14: y = 16'b0010001100000000;
        15: y = 16'b0010010100101111;
        16: y = 16'b0010011101001110;
        17: y = 16'b0010100101011100;
        18: y = 16'b0010101101010111;
        19: y = 16'b0010110101000000;
        20: y = 16'b0010111100010101;
        21: y = 16'b0011000011010101;
        22: y = 16'b0011001010000000;
        23: y = 16'b0011010000010100;
        24: y = 16'b0011010110010010;
        25: y = 16'b0011011011111001;
        26: y = 16'b0011100001001000;
        27: y = 16'b0011100101111101;
        28: y = 16'b0011101010011010;
        29: y = 16'b0011101110011101;
        30: y = 16'b0011110010000110;
        31: y = 16'b0011110101010101;
        32: y = 16'b0011111000001001;
        33: y = 16'b0011111010100001;
        34: y = 16'b0011111100011111;
        35: y = 16'b0011111110000000;
        36: y = 16'b0011111111000110;
        37: y = 16'b0011111111110000;
        38: y = 16'b0011111111111110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=369.99Hz, Fs=52734Hz, 16-bit, Volume 14/15 bit

module table_52734_Fs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 36;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001011001011;
        2: y = 16'b0000010110010100;
        3: y = 16'b0000100001011010;
        4: y = 16'b0000101100011101;
        5: y = 16'b0000110111011010;
        6: y = 16'b0001000010010000;
        7: y = 16'b0001001100111110;
        8: y = 16'b0001010111100011;
        9: y = 16'b0001100001111101;
        10: y = 16'b0001101100001011;
        11: y = 16'b0001110110001100;
        12: y = 16'b0001111111111111;
        13: y = 16'b0010001001100010;
        14: y = 16'b0010010010110100;
        15: y = 16'b0010011011110101;
        16: y = 16'b0010100100100010;
        17: y = 16'b0010101100111100;
        18: y = 16'b0010110101000000;
        19: y = 16'b0010111100101110;
        20: y = 16'b0011000100000101;
        21: y = 16'b0011001011000101;
        22: y = 16'b0011010001101011;
        23: y = 16'b0011010111111000;
        24: y = 16'b0011011101101011;
        25: y = 16'b0011100011000011;
        26: y = 16'b0011100111111111;
        27: y = 16'b0011101100011111;
        28: y = 16'b0011110000100010;
        29: y = 16'b0011110100001000;
        30: y = 16'b0011110111010000;
        31: y = 16'b0011111001111010;
        32: y = 16'b0011111100000101;
        33: y = 16'b0011111101110010;
        34: y = 16'b0011111111000000;
        35: y = 16'b0011111111101110;
        36: y = 16'b0011111111111110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=392.0Hz, Fs=52734Hz, 16-bit, Volume 14/15 bit

module table_52734_G
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 34;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001011110101;
        2: y = 16'b0000010111101000;
        3: y = 16'b0000100011010111;
        4: y = 16'b0000101111000010;
        5: y = 16'b0000111010100111;
        6: y = 16'b0001000110000011;
        7: y = 16'b0001010001010110;
        8: y = 16'b0001011100011110;
        9: y = 16'b0001100111011001;
        10: y = 16'b0001110010000110;
        11: y = 16'b0001111100100100;
        12: y = 16'b0010000110110000;
        13: y = 16'b0010010000101010;
        14: y = 16'b0010011010010000;
        15: y = 16'b0010100011100010;
        16: y = 16'b0010101100011100;
        17: y = 16'b0010110101000000;
        18: y = 16'b0010111101001010;
        19: y = 16'b0011000100111011;
        20: y = 16'b0011001100010001;
        21: y = 16'b0011010011001011;
        22: y = 16'b0011011001101000;
        23: y = 16'b0011011111101000;
        24: y = 16'b0011100101001001;
        25: y = 16'b0011101010001010;
        26: y = 16'b0011101110101100;
        27: y = 16'b0011110010101101;
        28: y = 16'b0011110110001101;
        29: y = 16'b0011111001001011;
        30: y = 16'b0011111011100111;
        31: y = 16'b0011111101100001;
        32: y = 16'b0011111110111000;
        33: y = 16'b0011111111101101;
        34: y = 16'b0011111111111110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=415.3Hz, Fs=52734Hz, 16-bit, Volume 14/15 bit

module table_52734_Gs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 32;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001100100100;
        2: y = 16'b0000011001000110;
        3: y = 16'b0000100101100100;
        4: y = 16'b0000110001111100;
        5: y = 16'b0000111110001101;
        6: y = 16'b0001001010010011;
        7: y = 16'b0001010110001111;
        8: y = 16'b0001100001111101;
        9: y = 16'b0001101101011100;
        10: y = 16'b0001111000101010;
        11: y = 16'b0010000011100110;
        12: y = 16'b0010001110001101;
        13: y = 16'b0010011000011111;
        14: y = 16'b0010100010011001;
        15: y = 16'b0010101011111001;
        16: y = 16'b0010110101000000;
        17: y = 16'b0010111101101010;
        18: y = 16'b0011000101110111;
        19: y = 16'b0011001101100110;
        20: y = 16'b0011010100110101;
        21: y = 16'b0011011011100011;
        22: y = 16'b0011100001110000;
        23: y = 16'b0011100111011001;
        24: y = 16'b0011101100011111;
        25: y = 16'b0011110001000000;
        26: y = 16'b0011110100111101;
        27: y = 16'b0011111000010011;
        28: y = 16'b0011111011000011;
        29: y = 16'b0011111101001101;
        30: y = 16'b0011111110101111;
        31: y = 16'b0011111111101010;
        32: y = 16'b0011111111111110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=440.0Hz, Fs=52734Hz, 16-bit, Volume 14/15 bit

module table_52734_A
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 30;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001101011001;
        2: y = 16'b0000011010110000;
        3: y = 16'b0000101000000011;
        4: y = 16'b0000110101001110;
        5: y = 16'b0001000010010000;
        6: y = 16'b0001001111000110;
        7: y = 16'b0001011011101111;
        8: y = 16'b0001101000000111;
        9: y = 16'b0001110100001101;
        10: y = 16'b0001111111111111;
        11: y = 16'b0010001011011010;
        12: y = 16'b0010010110011101;
        13: y = 16'b0010100001000110;
        14: y = 16'b0010101011010010;
        15: y = 16'b0010110101000000;
        16: y = 16'b0010111110001110;
        17: y = 16'b0011000110111011;
        18: y = 16'b0011001111000101;
        19: y = 16'b0011010110101011;
        20: y = 16'b0011011101101011;
        21: y = 16'b0011100100000100;
        22: y = 16'b0011101001110110;
        23: y = 16'b0011101110111110;
        24: y = 16'b0011110011011100;
        25: y = 16'b0011110111010000;
        26: y = 16'b0011111010011000;
        27: y = 16'b0011111100110100;
        28: y = 16'b0011111110100100;
        29: y = 16'b0011111111101000;
        30: y = 16'b0011111111111110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=466.16Hz, Fs=52734Hz, 16-bit, Volume 14/15 bit

module table_52734_As
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 28;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001110010111;
        2: y = 16'b0000011100101010;
        3: y = 16'b0000101010111000;
        4: y = 16'b0000111000111101;
        5: y = 16'b0001000110110111;
        6: y = 16'b0001010100100011;
        7: y = 16'b0001100001111101;
        8: y = 16'b0001101111000100;
        9: y = 16'b0001111011110100;
        10: y = 16'b0010001000001100;
        11: y = 16'b0010010100001000;
        12: y = 16'b0010011111100110;
        13: y = 16'b0010101010100100;
        14: y = 16'b0010110101000000;
        15: y = 16'b0010111110110111;
        16: y = 16'b0011001000001000;
        17: y = 16'b0011010000110001;
        18: y = 16'b0011011000101111;
        19: y = 16'b0011100000000010;
        20: y = 16'b0011100110101000;
        21: y = 16'b0011101100011111;
        22: y = 16'b0011110001100111;
        23: y = 16'b0011110101111110;
        24: y = 16'b0011111001100011;
        25: y = 16'b0011111100010111;
        26: y = 16'b0011111110010111;
        27: y = 16'b0011111111100100;
        28: y = 16'b0011111111111110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin((1/4)*2*pi*t*(F/Fs)), F=493.88Hz, Fs=52734Hz, 16-bit, Volume 14/15 bit

module table_52734_B
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 27;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001110111001;
        2: y = 16'b0000011101101110;
        3: y = 16'b0000101100011101;
        4: y = 16'b0000111011000010;
        5: y = 16'b0001001001011010;
        6: y = 16'b0001010111100011;
        7: y = 16'b0001100101011001;
        8: y = 16'b0001110010111000;
        9: y = 16'b0001111111111111;
        10: y = 16'b0010001100101010;
        11: y = 16'b0010011000110111;
        12: y = 16'b0010100100100010;
        13: y = 16'b0010101111101010;
        14: y = 16'b0010111010001100;
        15: y = 16'b0011000100000101;
        16: y = 16'b0011001101010100;
        17: y = 16'b0011010101110111;
        18: y = 16'b0011011101101011;
        19: y = 16'b0011100100101111;
        20: y = 16'b0011101011000010;
        21: y = 16'b0011110000100010;
        22: y = 16'b0011110101001110;
        23: y = 16'b0011111001000100;
        24: y = 16'b0011111100000101;
        25: y = 16'b0011111110001111;
        26: y = 16'b0011111111100010;
        27: y = 16'b0011111111111110;
        default: y = 16'b0;
        endcase

endmodule

