
module instruction_ram
#(
    parameter SIZE = 256
)
(
    input logic         clk,

    input  logic        mem_valid,
    output logic        mem_ready,

    input  logic [31:0] mem_addr,
    input  logic [3:0]  mem_wstrb,

    output logic [31:0] mem_rdata,
    input  logic [31:0] mem_wdata
);
    logic [31:0] memory [0:SIZE - 1];

    initial $readmemh ("program.hex", memory);

    always @(posedge clk) begin
		if (mem_valid) begin
			if (mem_addr < 1024) begin
				mem_rdata <= memory[mem_addr >> 2];
				if (mem_wstrb[0]) memory[mem_addr >> 2][ 7: 0] <= mem_wdata[ 7: 0];
				if (mem_wstrb[1]) memory[mem_addr >> 2][15: 8] <= mem_wdata[15: 8];
				if (mem_wstrb[2]) memory[mem_addr >> 2][23:16] <= mem_wdata[23:16];
				if (mem_wstrb[3]) memory[mem_addr >> 2][31:24] <= mem_wdata[31:24];
			end
		end
	end

    assign mem_ready = 1'b1;

endmodule
