`include "../omdazz_epm570/board_specific_top.sv"
