`define USE_HUB75E_LED_MATRIX_64x64
`include "../tang_primer_25k_pmod_vga/board_specific_top.sv"
