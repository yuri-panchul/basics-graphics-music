`include "config.svh"

module lab_top
# (
    parameter  clk_mhz       = 50,
               w_key         = 4,
               w_sw          = 8,
               w_led         = 8,
               w_digit       = 8,
               w_gpio        = 100,

               screen_width  = 640,
               screen_height = 480,

               w_red         = 4,
               w_green       = 4,
               w_blue        = 4,

               w_x           = $clog2 ( screen_width  ),
               w_y           = $clog2 ( screen_height )
)
(
    input                        clk,
    input                        slow_clk,
    input                        rst,

    // Keys, switches, LEDs

    input        [w_key   - 1:0] key,
    input        [w_sw    - 1:0] sw,
    output logic [w_led   - 1:0] led,

    // A dynamic seven-segment display

    output logic [          7:0] abcdefgh,
    output logic [w_digit - 1:0] digit,

    // Graphics

    input        [w_x     - 1:0] x,
    input        [w_y     - 1:0] y,

    output logic [w_red   - 1:0] red,
    output logic [w_green - 1:0] green,
    output logic [w_blue  - 1:0] blue,

    // Microphone, sound output and UART

    input        [         23:0] mic,
    output       [         15:0] sound,

    input                        uart_rx,
    output                       uart_tx,

    // General-purpose Input/Output

    inout        [w_gpio  - 1:0] gpio
);

    //------------------------------------------------------------------------

    // assign led        = '0;
       assign abcdefgh   = '0;
       assign digit      = '0;
       assign red        = '0;
       assign green      = '0;
       assign blue       = '0;
       assign sound      = '0;
       assign uart_tx    = '1;

    //------------------------------------------------------------------------

    localparam w_in = 8;
    wire [w_in - 1:0] in;

    generate
        if (w_key < w_in && w_sw >= w_in)
        begin : use_switches
            assign in = w_in' (sw);
        end
        else
        begin : use_keys
            assign in = w_in' (key);
        end
    endgenerate

    //------------------------------------------------------------------------

    mux_2_1_using_conditional_operator mux_1
    (
        .a   ( in  [1]   ),
        .b   ( in  [0]   ),
        .sel ( in  [2]   ),
        .out ( led [0]   )
    );

    mux_2_1_using_gates mux_2
    (
        .a   ( in  [1]   ),
        .b   ( in  [0]   ),
        .sel ( in  [2]   ),
        .out ( led [1]   )
    );

    mux_2_1_width_3_using_if mux_3
    (
        .a   ( in  [5:3] ),
        .b   ( in  [2:0] ),
        .sel ( in  [7]   ),
        .out ( led [7:5] )
    );

    mux_5_1_using_case mux_4
    (
        .a   ( in  [4]   ),
        .b   ( in  [3]   ),
        .c   ( in  [2]   ),
        .d   ( in  [1]   ),
        .e   ( in  [0]   ),
        .sel ( in  [7:5] ),
        .out ( led [2]   )
    );

    mux_4_1_using_indexing mux_5
    (
        .in  ( in  [3:0] ),
        .sel ( in  [7:6] ),
        .out ( led [3]   )
    );

endmodule
