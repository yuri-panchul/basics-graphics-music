`define USE_PMOD_DVI
`include "../tang_primer_25k_pmod_vga/board_specific_top.sv"
