`include "config.svh"

module tb;

  localparam clk_mhz = 1,
             w_key   = 4,
             w_sw    = 8,
             w_led   = 8,
             w_digit = 8,
             w_gpio  = 20;

  //--------------------------------------------------------------------------

  logic       clk;
  logic       rst;
  logic [3:0] key;
  logic [7:0] sw;

  //--------------------------------------------------------------------------

  top
  # (
    .clk_mhz ( clk_mhz ),
    .w_key   ( w_key   ),
    .w_sw    ( w_sw    ),
    .w_led   ( w_led   ),
    .w_digit ( w_digit ),
    .w_gpio  ( w_gpio  )
  )
  i_top
  (
    .clk ( clk ),
    .rst ( rst ),
    .key ( key ),
    .sw  ( sw  )
  );

  //--------------------------------------------------------------------------

  initial
  begin
    `ifdef __ICARUS__
      $dumpvars;
    `endif

    repeat (8)
    begin
       #10
       key <= $urandom ();
       sw  <= $urandom ();
    end

    $finish;
  end

endmodule
