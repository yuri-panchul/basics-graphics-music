module sine_table(
    input  logic [7:0] idx_i,
    output logic [7:0] sine_o 
);

    always_comb begin
        case(idx_i)
           8'd0 : sine_o = 8'h00;
           8'd1 : sine_o = 8'h00;
           8'd2 : sine_o = 8'h00;
           8'd3 : sine_o = 8'h00;
           8'd4 : sine_o = 8'h00;
           8'd5 : sine_o = 8'h00;
           8'd6 : sine_o = 8'h00;
           8'd7 : sine_o = 8'h00;
           8'd8 : sine_o = 8'h01;
           8'd9 : sine_o = 8'h01;
           8'd10 : sine_o = 8'h01;
           8'd11 : sine_o = 8'h01;
           8'd12 : sine_o = 8'h01;
           8'd13 : sine_o = 8'h02;
           8'd14 : sine_o = 8'h02;
           8'd15 : sine_o = 8'h02;
           8'd16 : sine_o = 8'h02;
           8'd17 : sine_o = 8'h03;
           8'd18 : sine_o = 8'h03;
           8'd19 : sine_o = 8'h03;
           8'd20 : sine_o = 8'h04;
           8'd21 : sine_o = 8'h04;
           8'd22 : sine_o = 8'h05;
           8'd23 : sine_o = 8'h05;
           8'd24 : sine_o = 8'h06;
           8'd25 : sine_o = 8'h06;
           8'd26 : sine_o = 8'h06;
           8'd27 : sine_o = 8'h07;
           8'd28 : sine_o = 8'h08;
           8'd29 : sine_o = 8'h08;
           8'd30 : sine_o = 8'h09;
           8'd31 : sine_o = 8'h09;
           8'd32 : sine_o = 8'h0A;
           8'd33 : sine_o = 8'h0A;
           8'd34 : sine_o = 8'h0B;
           8'd35 : sine_o = 8'h0C;
           8'd36 : sine_o = 8'h0C;
           8'd37 : sine_o = 8'h0D;
           8'd38 : sine_o = 8'h0E;
           8'd39 : sine_o = 8'h0E;
           8'd40 : sine_o = 8'h0F;
           8'd41 : sine_o = 8'h10;
           8'd42 : sine_o = 8'h11;
           8'd43 : sine_o = 8'h11;
           8'd44 : sine_o = 8'h12;
           8'd45 : sine_o = 8'h13;
           8'd46 : sine_o = 8'h14;
           8'd47 : sine_o = 8'h15;
           8'd48 : sine_o = 8'h16;
           8'd49 : sine_o = 8'h17;
           8'd50 : sine_o = 8'h17;
           8'd51 : sine_o = 8'h18;
           8'd52 : sine_o = 8'h19;
           8'd53 : sine_o = 8'h1A;
           8'd54 : sine_o = 8'h1B;
           8'd55 : sine_o = 8'h1C;
           8'd56 : sine_o = 8'h1D;
           8'd57 : sine_o = 8'h1E;
           8'd58 : sine_o = 8'h1F;
           8'd59 : sine_o = 8'h20;
           8'd60 : sine_o = 8'h21;
           8'd61 : sine_o = 8'h22;
           8'd62 : sine_o = 8'h23;
           8'd63 : sine_o = 8'h25;
           8'd64 : sine_o = 8'h26;
           8'd65 : sine_o = 8'h27;
           8'd66 : sine_o = 8'h28;
           8'd67 : sine_o = 8'h29;
           8'd68 : sine_o = 8'h2A;
           8'd69 : sine_o = 8'h2B;
           8'd70 : sine_o = 8'h2D;
           8'd71 : sine_o = 8'h2E;
           8'd72 : sine_o = 8'h2F;
           8'd73 : sine_o = 8'h30;
           8'd74 : sine_o = 8'h31;
           8'd75 : sine_o = 8'h33;
           8'd76 : sine_o = 8'h34;
           8'd77 : sine_o = 8'h35;
           8'd78 : sine_o = 8'h36;
           8'd79 : sine_o = 8'h38;
           8'd80 : sine_o = 8'h39;
           8'd81 : sine_o = 8'h3A;
           8'd82 : sine_o = 8'h3C;
           8'd83 : sine_o = 8'h3D;
           8'd84 : sine_o = 8'h3E;
           8'd85 : sine_o = 8'h40;
           8'd86 : sine_o = 8'h41;
           8'd87 : sine_o = 8'h42;
           8'd88 : sine_o = 8'h44;
           8'd89 : sine_o = 8'h45;
           8'd90 : sine_o = 8'h47;
           8'd91 : sine_o = 8'h48;
           8'd92 : sine_o = 8'h49;
           8'd93 : sine_o = 8'h4B;
           8'd94 : sine_o = 8'h4C;
           8'd95 : sine_o = 8'h4E;
           8'd96 : sine_o = 8'h4F;
           8'd97 : sine_o = 8'h51;
           8'd98 : sine_o = 8'h52;
           8'd99 : sine_o = 8'h54;
           8'd100 : sine_o = 8'h55;
           8'd101 : sine_o = 8'h57;
           8'd102 : sine_o = 8'h58;
           8'd103 : sine_o = 8'h5A;
           8'd104 : sine_o = 8'h5B;
           8'd105 : sine_o = 8'h5D;
           8'd106 : sine_o = 8'h5E;
           8'd107 : sine_o = 8'h60;
           8'd108 : sine_o = 8'h61;
           8'd109 : sine_o = 8'h63;
           8'd110 : sine_o = 8'h64;
           8'd111 : sine_o = 8'h66;
           8'd112 : sine_o = 8'h67;
           8'd113 : sine_o = 8'h69;
           8'd114 : sine_o = 8'h6A;
           8'd115 : sine_o = 8'h6C;
           8'd116 : sine_o = 8'h6D;
           8'd117 : sine_o = 8'h6F;
           8'd118 : sine_o = 8'h71;
           8'd119 : sine_o = 8'h72;
           8'd120 : sine_o = 8'h74;
           8'd121 : sine_o = 8'h75;
           8'd122 : sine_o = 8'h77;
           8'd123 : sine_o = 8'h78;
           8'd124 : sine_o = 8'h7A;
           8'd125 : sine_o = 8'h7C;
           8'd126 : sine_o = 8'h7D;
           8'd127 : sine_o = 8'h7F;
           8'd128 : sine_o = 8'h80;
           8'd129 : sine_o = 8'h82;
           8'd130 : sine_o = 8'h83;
           8'd131 : sine_o = 8'h85;
           8'd132 : sine_o = 8'h87;
           8'd133 : sine_o = 8'h88;
           8'd134 : sine_o = 8'h8A;
           8'd135 : sine_o = 8'h8B;
           8'd136 : sine_o = 8'h8D;
           8'd137 : sine_o = 8'h8E;
           8'd138 : sine_o = 8'h90;
           8'd139 : sine_o = 8'h92;
           8'd140 : sine_o = 8'h93;
           8'd141 : sine_o = 8'h95;
           8'd142 : sine_o = 8'h96;
           8'd143 : sine_o = 8'h98;
           8'd144 : sine_o = 8'h99;
           8'd145 : sine_o = 8'h9B;
           8'd146 : sine_o = 8'h9C;
           8'd147 : sine_o = 8'h9E;
           8'd148 : sine_o = 8'h9F;
           8'd149 : sine_o = 8'hA1;
           8'd150 : sine_o = 8'hA2;
           8'd151 : sine_o = 8'hA4;
           8'd152 : sine_o = 8'hA5;
           8'd153 : sine_o = 8'hA7;
           8'd154 : sine_o = 8'hA8;
           8'd155 : sine_o = 8'hAA;
           8'd156 : sine_o = 8'hAB;
           8'd157 : sine_o = 8'hAD;
           8'd158 : sine_o = 8'hAE;
           8'd159 : sine_o = 8'hB0;
           8'd160 : sine_o = 8'hB1;
           8'd161 : sine_o = 8'hB3;
           8'd162 : sine_o = 8'hB4;
           8'd163 : sine_o = 8'hB6;
           8'd164 : sine_o = 8'hB7;
           8'd165 : sine_o = 8'hB8;
           8'd166 : sine_o = 8'hBA;
           8'd167 : sine_o = 8'hBB;
           8'd168 : sine_o = 8'hBD;
           8'd169 : sine_o = 8'hBE;
           8'd170 : sine_o = 8'hBF;
           8'd171 : sine_o = 8'hC1;
           8'd172 : sine_o = 8'hC2;
           8'd173 : sine_o = 8'hC3;
           8'd174 : sine_o = 8'hC5;
           8'd175 : sine_o = 8'hC6;
           8'd176 : sine_o = 8'hC7;
           8'd177 : sine_o = 8'hC9;
           8'd178 : sine_o = 8'hCA;
           8'd179 : sine_o = 8'hCB;
           8'd180 : sine_o = 8'hCC;
           8'd181 : sine_o = 8'hCE;
           8'd182 : sine_o = 8'hCF;
           8'd183 : sine_o = 8'hD0;
           8'd184 : sine_o = 8'hD1;
           8'd185 : sine_o = 8'hD2;
           8'd186 : sine_o = 8'hD4;
           8'd187 : sine_o = 8'hD5;
           8'd188 : sine_o = 8'hD6;
           8'd189 : sine_o = 8'hD7;
           8'd190 : sine_o = 8'hD8;
           8'd191 : sine_o = 8'hD9;
           8'd192 : sine_o = 8'hDA;
           8'd193 : sine_o = 8'hDC;
           8'd194 : sine_o = 8'hDD;
           8'd195 : sine_o = 8'hDE;
           8'd196 : sine_o = 8'hDF;
           8'd197 : sine_o = 8'hE0;
           8'd198 : sine_o = 8'hE1;
           8'd199 : sine_o = 8'hE2;
           8'd200 : sine_o = 8'hE3;
           8'd201 : sine_o = 8'hE4;
           8'd202 : sine_o = 8'hE5;
           8'd203 : sine_o = 8'hE6;
           8'd204 : sine_o = 8'hE7;
           8'd205 : sine_o = 8'hE8;
           8'd206 : sine_o = 8'hE8;
           8'd207 : sine_o = 8'hE9;
           8'd208 : sine_o = 8'hEA;
           8'd209 : sine_o = 8'hEB;
           8'd210 : sine_o = 8'hEC;
           8'd211 : sine_o = 8'hED;
           8'd212 : sine_o = 8'hEE;
           8'd213 : sine_o = 8'hEE;
           8'd214 : sine_o = 8'hEF;
           8'd215 : sine_o = 8'hF0;
           8'd216 : sine_o = 8'hF1;
           8'd217 : sine_o = 8'hF1;
           8'd218 : sine_o = 8'hF2;
           8'd219 : sine_o = 8'hF3;
           8'd220 : sine_o = 8'hF3;
           8'd221 : sine_o = 8'hF4;
           8'd222 : sine_o = 8'hF5;
           8'd223 : sine_o = 8'hF5;
           8'd224 : sine_o = 8'hF6;
           8'd225 : sine_o = 8'hF6;
           8'd226 : sine_o = 8'hF7;
           8'd227 : sine_o = 8'hF7;
           8'd228 : sine_o = 8'hF8;
           8'd229 : sine_o = 8'hF9;
           8'd230 : sine_o = 8'hF9;
           8'd231 : sine_o = 8'hF9;
           8'd232 : sine_o = 8'hFA;
           8'd233 : sine_o = 8'hFA;
           8'd234 : sine_o = 8'hFB;
           8'd235 : sine_o = 8'hFB;
           8'd236 : sine_o = 8'hFC;
           8'd237 : sine_o = 8'hFC;
           8'd238 : sine_o = 8'hFC;
           8'd239 : sine_o = 8'hFD;
           8'd240 : sine_o = 8'hFD;
           8'd241 : sine_o = 8'hFD;
           8'd242 : sine_o = 8'hFD;
           8'd243 : sine_o = 8'hFE;
           8'd244 : sine_o = 8'hFE;
           8'd245 : sine_o = 8'hFE;
           8'd246 : sine_o = 8'hFE;
           8'd247 : sine_o = 8'hFE;
           8'd248 : sine_o = 8'hFF;
           8'd249 : sine_o = 8'hFF;
           8'd250 : sine_o = 8'hFF;
           8'd251 : sine_o = 8'hFF;
           8'd252 : sine_o = 8'hFF;
           8'd253 : sine_o = 8'hFF;
           8'd254 : sine_o = 8'hFF;
           8'd255 : sine_o = 8'hFF;
        endcase        
    end    

endmodule