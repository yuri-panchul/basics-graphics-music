`include "config.svh"

module top
# (
  parameter clk_mhz = 50,
            w_key   = 4,
            w_sw    = 8,
            w_led   = 8,
            w_digit = 8,
            w_gpio  = 20
)
(
  input                        clk,
  input                        rst,

  // Keys, switches, LEDs

  input        [w_key   - 1:0] key,
  input        [w_sw    - 1:0] sw,
  output logic [w_led   - 1:0] led,

  // A dynamic seven-segment display

  output logic [          7:0] abcdefgh,
  output logic [w_digit - 1:0] digit,

  // VGA

  output logic                 vsync,
  output logic                 hsync,
  output logic [          3:0] red,
  output logic [          3:0] green,
  output logic [          3:0] blue,

  // General-purpose Input/Output

  inout  logic [w_gpio  - 1:0] gpio
);

  //--------------------------------------------------------------------------

  // assign led      = '0;
  // assign abcdefgh = '0;
  // assign digit    = '0;
     assign vsync    = '0;
     assign hsync    = '0;
     assign red      = '0;
     assign green    = '0;
     assign blue     = '0;

  //--------------------------------------------------------------------------

  // Exercise 1: Free running counter.
  // How do you change the speed of LED blinking?
  // Try different bit slices to display.

  logic [31:0] cnt;

  always_ff @ (posedge clk or posedge rst)
    if (rst)
      cnt <= '0;
    else
      cnt <= cnt + 1'd1;

  assign led      = cnt [ $left ( led      ) -: w_led   ];
  assign abcdefgh = cnt [ $left ( abcdefgh ) -: 8       ];
  assign digit    = cnt [ $left ( digit    ) -: w_digit ];

  // Exercise 2: Key-controlled counter.
  // Comment out the code above.
  // Uncomment and synthesize the code below.
  // Press the key to see the counter incrementing.
  //
  // Change the design, for example:
  //
  // 1. One key is used to increment, another to decrement.
  //
  // 2. Two counters controlled by different keys
  // displayed in different groups of LEDs.

  /*

  wire any_key = | key;

  logic any_key_r;

  always_ff @ (posedge clk or posedge rst)
    if (rst)
      any_key_r <= '0;
    else
      any_key_r <= any_key;

  wire any_key_pressed = ~ any_key & any_key_r;

  logic [3:0] cnt;

  always_ff @ (posedge clk or posedge rst)
    if (rst)
      cnt <= '0;
    else if (any_key_pressed)
      cnt <= cnt + 1'd1;

  */

endmodule
