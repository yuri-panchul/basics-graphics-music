`include "../omdazz/board_specific_top.sv"
