`ifndef LAB_SPECIFIC_CONFIG_SVH
`define LAB_SPECIFIC_CONFIG_SVH

// The following setting is needed for Gowin boards
   `define INSTANTIATE_TM1638_BOARD_CONTROLLER_MODULE

// HCW-132 variant of LED & KEY TM1638 board controller
// `define USE_HCW132_VARIANT_OF_TM1638_BOARD_CONTROLLER_MODULE

// `define EMULATE_DYNAMIC_7SEG_ON_STATIC_WITHOUT_STICKY_FLOPS

// `define DUPLICATE_TM1638_SIGNALS_WITH_REGULAR
// `define CONCAT_REGULAR_SIGNALS_AND_TM
   `define CONCAT_TM1638_SIGNALS_AND_REGULAR

`endif  // `ifndef LAB_SPECIFIC_CONFIG_SVH
