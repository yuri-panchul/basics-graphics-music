`include "../nexys_a7/board_specific_top.sv"
