// This module is created based on https://github.com/sipeed/TangNano-9K-example/lcd_led/src/VGAMod.v
// Timining were take from https://github.com/HASwitchPlate/openHASP/blob/master/user_setups/esp32s3/sunton-esp32-s3-tft.ini

module lcd_480_272_ml6485
(
    input                   nRST,

    input                   PixelClk,

    output                  LCD_DE,
    output                  LCD_HSYNC,
    output                  LCD_VSYNC,

    // Modified for basic-graphics-music: Removed LCD_RGB ports.
    // These output signals are assigned in the top module code
    // using input from lab_top module.

    /*
    output          [4:0]   LCD_B,
    output          [5:0]   LCD_G,
    output          [4:0]   LCD_R
    */

    // Modified for basic-graphics-music: Added x and y outputs

    output [9:0] x,
    output [8:0] y
);

    reg         [15:0]  PixelCount;
    reg         [15:0]  LineCount;

    localparam      V_BackPorch = 16'd12;
    localparam      V_Pluse     = 16'd4;
    localparam      HightPixel  = 16'd272;
    localparam      V_FrontPorch= 16'd64;

    localparam      H_BackPorch = 16'd43;
    localparam      H_Pluse     = 16'd4;
    localparam      WidthPixel  = 16'd480;
    localparam      H_FrontPorch= 16'd64;

    parameter       BarCount    = 16; // RGB565
    localparam      Width_bar   = WidthPixel / 16;

    localparam      PixelForHS  =   WidthPixel + H_BackPorch + H_FrontPorch;
    localparam      LineForVS   =   HightPixel + V_BackPorch + V_FrontPorch;

    always @(  posedge PixelClk or negedge nRST  )begin
        if( !nRST ) begin
            LineCount       <=  16'b0;
            PixelCount      <=  16'b0;
            end
        else if(  PixelCount  ==  PixelForHS ) begin
            PixelCount      <=  16'b0;
            LineCount       <=  LineCount + 1'b1;
            end
        else if(  LineCount  == LineForVS  ) begin
            LineCount       <=  16'b0;
            PixelCount      <=  16'b0;
            end
        else
            PixelCount      <=  PixelCount + 1'b1;
    end

    reg            [9:0]  Data_R;
    reg            [9:0]  Data_G;
    reg            [9:0]  Data_B;

    always @(  posedge PixelClk or negedge nRST  )begin
        if( !nRST ) begin
            Data_R <= 9'b0;
            Data_G <= 9'b0;
            Data_B <= 9'b0;
            end
    end
    //注意这里HSYNC和VSYNC负极性
    assign  LCD_HSYNC = (( PixelCount >= H_Pluse)&&( PixelCount <= (PixelForHS-H_FrontPorch))) ? 1'b0 : 1'b1;
    //assign  LCD_VSYNC = ((( LineCount  >= 0 )&&( LineCount  <= (V_Pluse-1) )) ) ? 1'b1 : 1'b0;        //这里不减一的话，图片底部会往下拖尾？
    assign  LCD_VSYNC = ((( LineCount  >= V_Pluse )&&( LineCount  <= (LineForVS-0) )) ) ? 1'b0 : 1'b1;
    //assign  FIFO_RST  = (( PixelCount ==0)) ? 1'b1 : 1'b0;  //留给主机H_BackPorch的时间进入中断，发送数据

    assign  LCD_DE = (  ( PixelCount >= H_BackPorch )&&
                        ( PixelCount <= PixelForHS-H_FrontPorch ) &&
                        ( LineCount >= V_BackPorch ) &&
                        ( LineCount <= LineForVS-V_FrontPorch-1 ))  ? 1'b1 : 1'b0;
                        //这里不减一，会抖动

    // Modified for basic-graphics-music: Removed LCD_RGB port assignments.
    // These output signals are assigned in the top module code
    // using input from lab_top module.

    `ifdef COMMENTED_OUT

    // assign  LCD_R   =   (PixelCount<200)? 5'b00000 :
    //                     (PixelCount<240 ? 5'b00001 :
    //                     (PixelCount<280 ? 5'b00010 :
    //                     (PixelCount<320 ? 5'b00100 :
    //                     (PixelCount<360 ? 5'b01000 :
    //                     (PixelCount<400 ? 5'b10000 :  5'b00000 )))));

    // assign  LCD_G   =   (PixelCount<400)? 6'b000000 :
    //                     (PixelCount<440 ? 6'b000001 :
    //                     (PixelCount<480 ? 6'b000010 :
    //                     (PixelCount<520 ? 6'b000100 :
    //                     (PixelCount<560 ? 6'b001000 :
    //                     (PixelCount<600 ? 6'b010000 :
    //                     (PixelCount<640 ? 6'b100000 : 6'b000000 ))))));

    // assign  LCD_B   =   (PixelCount<640)? 5'b00000 :
    //                     (PixelCount<680 ? 5'b00001 :
    //                     (PixelCount<720 ? 5'b00010 :
    //                     (PixelCount<760 ? 5'b00100 :
    //                     (PixelCount<800 ? 5'b01000 :
    //                     (PixelCount<840 ? 5'b10000 :  5'b00000 )))));

    assign  LCD_R   =   PixelCount < H_BackPorch + Width_bar *  0    ? 5'b00000 :
                        PixelCount < H_BackPorch + Width_bar *  1    ? 5'b00001 :
                        PixelCount < H_BackPorch + Width_bar *  2    ? 5'b00010 :
                        PixelCount < H_BackPorch + Width_bar *  3    ? 5'b00100 :
                        PixelCount < H_BackPorch + Width_bar *  4    ? 5'b01000 :
                        PixelCount < H_BackPorch + Width_bar *  5    ? 5'b10000 :  5'b00000 ;

    assign  LCD_G   =   PixelCount < H_BackPorch + Width_bar *  6    ? 6'b000001 :
                        PixelCount < H_BackPorch + Width_bar *  7    ? 6'b000010 :
                        PixelCount < H_BackPorch + Width_bar *  8    ? 6'b000100 :
                        PixelCount < H_BackPorch + Width_bar *  9    ? 6'b001000 :
                        PixelCount < H_BackPorch + Width_bar *  10   ? 6'b010000 :
                        PixelCount < H_BackPorch + Width_bar *  11   ? 6'b100000 : 6'b000000 ;

    assign  LCD_B   =   PixelCount < H_BackPorch + Width_bar *  12   ? 5'b00001 :
                        PixelCount < H_BackPorch + Width_bar *  13   ? 5'b00010 :
                        PixelCount < H_BackPorch + Width_bar *  14   ? 5'b00100 :
                        PixelCount < H_BackPorch + Width_bar *  15   ? 5'b01000 :
                        PixelCount < H_BackPorch + Width_bar *  16   ? 5'b10000 :  5'b00000 ;

    `endif

    // Modified for basic-graphics-music: Added x and y outputs

    assign x = 10' (PixelCount - H_BackPorch);
    assign y =  9' (LineCount  - V_BackPorch);

endmodule
