`define FORCE_NO_INSTANTIATE_GRAPHICS_INTERFACE_MODULE
`include "../tang_primer_20k_dock_hdmi_tm1638/board_specific_top.sv"
