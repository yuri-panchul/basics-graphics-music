`define  COMPENSATE_DEFECTIVE_BOARD_WITH_DIGIT_0_NOT_WORKING
`include "../zeowaa/board_specific_top.sv"
