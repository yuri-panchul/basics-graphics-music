// y(t) = sin(2*pi*F*t), F=261.63Hz, Fs=96000Hz, 16-bit

module lut_C
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 365;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001000110010;
        2: y = 16'b0000010001100101;
        3: y = 16'b0000011010010111;
        4: y = 16'b0000100011001000;
        5: y = 16'b0000101011111001;
        6: y = 16'b0000110100101001;
        7: y = 16'b0000111101011000;
        8: y = 16'b0001000110000110;
        9: y = 16'b0001001110110011;
        10: y = 16'b0001010111011110;
        11: y = 16'b0001100000000111;
        12: y = 16'b0001101000101111;
        13: y = 16'b0001110001010100;
        14: y = 16'b0001111001111000;
        15: y = 16'b0010000010011001;
        16: y = 16'b0010001010111000;
        17: y = 16'b0010010011010100;
        18: y = 16'b0010011011101101;
        19: y = 16'b0010100100000011;
        20: y = 16'b0010101100010111;
        21: y = 16'b0010110100100111;
        22: y = 16'b0010111100110011;
        23: y = 16'b0011000100111100;
        24: y = 16'b0011001101000010;
        25: y = 16'b0011010101000011;
        26: y = 16'b0011011101000001;
        27: y = 16'b0011100100111010;
        28: y = 16'b0011101100101111;
        29: y = 16'b0011110100011111;
        30: y = 16'b0011111100001011;
        31: y = 16'b0100000011110010;
        32: y = 16'b0100001011010101;
        33: y = 16'b0100010010110010;
        34: y = 16'b0100011010001010;
        35: y = 16'b0100100001011101;
        36: y = 16'b0100101000101010;
        37: y = 16'b0100101111110010;
        38: y = 16'b0100110110110011;
        39: y = 16'b0100111101110000;
        40: y = 16'b0101000100100110;
        41: y = 16'b0101001011010110;
        42: y = 16'b0101010001111111;
        43: y = 16'b0101011000100011;
        44: y = 16'b0101011110111111;
        45: y = 16'b0101100101010110;
        46: y = 16'b0101101011100101;
        47: y = 16'b0101110001101110;
        48: y = 16'b0101110111101111;
        49: y = 16'b0101111101101010;
        50: y = 16'b0110000011011101;
        51: y = 16'b0110001001001001;
        52: y = 16'b0110001110101110;
        53: y = 16'b0110010100001011;
        54: y = 16'b0110011001100000;
        55: y = 16'b0110011110101110;
        56: y = 16'b0110100011110100;
        57: y = 16'b0110101000110010;
        58: y = 16'b0110101101101000;
        59: y = 16'b0110110010010110;
        60: y = 16'b0110110110111100;
        61: y = 16'b0110111011011001;
        62: y = 16'b0110111111101110;
        63: y = 16'b0111000011111011;
        64: y = 16'b0111000111111111;
        65: y = 16'b0111001011111010;
        66: y = 16'b0111001111101101;
        67: y = 16'b0111010011010111;
        68: y = 16'b0111010110111000;
        69: y = 16'b0111011010010001;
        70: y = 16'b0111011101100000;
        71: y = 16'b0111100000100111;
        72: y = 16'b0111100011100100;
        73: y = 16'b0111100110011000;
        74: y = 16'b0111101001000011;
        75: y = 16'b0111101011100101;
        76: y = 16'b0111101101111110;
        77: y = 16'b0111110000001101;
        78: y = 16'b0111110010010011;
        79: y = 16'b0111110100001111;
        80: y = 16'b0111110110000011;
        81: y = 16'b0111110111101100;
        82: y = 16'b0111111001001100;
        83: y = 16'b0111111010100011;
        84: y = 16'b0111111011110000;
        85: y = 16'b0111111100110011;
        86: y = 16'b0111111101101101;
        87: y = 16'b0111111110011101;
        88: y = 16'b0111111111000100;
        89: y = 16'b0111111111100001;
        90: y = 16'b0111111111110100;
        91: y = 16'b0111111111111110;
        92: y = 16'b0111111111111110;
        93: y = 16'b0111111111110100;
        94: y = 16'b0111111111100001;
        95: y = 16'b0111111111000100;
        96: y = 16'b0111111110011101;
        97: y = 16'b0111111101101101;
        98: y = 16'b0111111100110011;
        99: y = 16'b0111111011110000;
        100: y = 16'b0111111010100011;
        101: y = 16'b0111111001001100;
        102: y = 16'b0111110111101100;
        103: y = 16'b0111110110000011;
        104: y = 16'b0111110100001111;
        105: y = 16'b0111110010010011;
        106: y = 16'b0111110000001101;
        107: y = 16'b0111101101111110;
        108: y = 16'b0111101011100101;
        109: y = 16'b0111101001000011;
        110: y = 16'b0111100110011000;
        111: y = 16'b0111100011100100;
        112: y = 16'b0111100000100111;
        113: y = 16'b0111011101100000;
        114: y = 16'b0111011010010001;
        115: y = 16'b0111010110111000;
        116: y = 16'b0111010011010111;
        117: y = 16'b0111001111101101;
        118: y = 16'b0111001011111010;
        119: y = 16'b0111000111111111;
        120: y = 16'b0111000011111011;
        121: y = 16'b0110111111101110;
        122: y = 16'b0110111011011001;
        123: y = 16'b0110110110111100;
        124: y = 16'b0110110010010110;
        125: y = 16'b0110101101101000;
        126: y = 16'b0110101000110010;
        127: y = 16'b0110100011110100;
        128: y = 16'b0110011110101110;
        129: y = 16'b0110011001100000;
        130: y = 16'b0110010100001011;
        131: y = 16'b0110001110101110;
        132: y = 16'b0110001001001001;
        133: y = 16'b0110000011011101;
        134: y = 16'b0101111101101010;
        135: y = 16'b0101110111101111;
        136: y = 16'b0101110001101110;
        137: y = 16'b0101101011100101;
        138: y = 16'b0101100101010110;
        139: y = 16'b0101011110111111;
        140: y = 16'b0101011000100011;
        141: y = 16'b0101010001111111;
        142: y = 16'b0101001011010110;
        143: y = 16'b0101000100100110;
        144: y = 16'b0100111101110000;
        145: y = 16'b0100110110110011;
        146: y = 16'b0100101111110010;
        147: y = 16'b0100101000101010;
        148: y = 16'b0100100001011101;
        149: y = 16'b0100011010001010;
        150: y = 16'b0100010010110010;
        151: y = 16'b0100001011010101;
        152: y = 16'b0100000011110010;
        153: y = 16'b0011111100001011;
        154: y = 16'b0011110100011111;
        155: y = 16'b0011101100101111;
        156: y = 16'b0011100100111010;
        157: y = 16'b0011011101000001;
        158: y = 16'b0011010101000011;
        159: y = 16'b0011001101000010;
        160: y = 16'b0011000100111100;
        161: y = 16'b0010111100110011;
        162: y = 16'b0010110100100111;
        163: y = 16'b0010101100010111;
        164: y = 16'b0010100100000011;
        165: y = 16'b0010011011101101;
        166: y = 16'b0010010011010100;
        167: y = 16'b0010001010111000;
        168: y = 16'b0010000010011001;
        169: y = 16'b0001111001111000;
        170: y = 16'b0001110001010100;
        171: y = 16'b0001101000101111;
        172: y = 16'b0001100000000111;
        173: y = 16'b0001010111011110;
        174: y = 16'b0001001110110011;
        175: y = 16'b0001000110000110;
        176: y = 16'b0000111101011000;
        177: y = 16'b0000110100101001;
        178: y = 16'b0000101011111001;
        179: y = 16'b0000100011001000;
        180: y = 16'b0000011010010111;
        181: y = 16'b0000010001100101;
        182: y = 16'b0000001000110010;
        183: y = 16'b0000000000000000;
        184: y = 16'b1111110111001110;
        185: y = 16'b1111101110011011;
        186: y = 16'b1111100101101001;
        187: y = 16'b1111011100111000;
        188: y = 16'b1111010100000111;
        189: y = 16'b1111001011010111;
        190: y = 16'b1111000010101000;
        191: y = 16'b1110111001111010;
        192: y = 16'b1110110001001101;
        193: y = 16'b1110101000100010;
        194: y = 16'b1110011111111001;
        195: y = 16'b1110010111010001;
        196: y = 16'b1110001110101100;
        197: y = 16'b1110000110001000;
        198: y = 16'b1101111101100111;
        199: y = 16'b1101110101001000;
        200: y = 16'b1101101100101100;
        201: y = 16'b1101100100010011;
        202: y = 16'b1101011011111101;
        203: y = 16'b1101010011101001;
        204: y = 16'b1101001011011001;
        205: y = 16'b1101000011001101;
        206: y = 16'b1100111011000100;
        207: y = 16'b1100110010111110;
        208: y = 16'b1100101010111101;
        209: y = 16'b1100100010111111;
        210: y = 16'b1100011011000110;
        211: y = 16'b1100010011010001;
        212: y = 16'b1100001011100001;
        213: y = 16'b1100000011110101;
        214: y = 16'b1011111100001110;
        215: y = 16'b1011110100101011;
        216: y = 16'b1011101101001110;
        217: y = 16'b1011100101110110;
        218: y = 16'b1011011110100011;
        219: y = 16'b1011010111010110;
        220: y = 16'b1011010000001110;
        221: y = 16'b1011001001001101;
        222: y = 16'b1011000010010000;
        223: y = 16'b1010111011011010;
        224: y = 16'b1010110100101010;
        225: y = 16'b1010101110000001;
        226: y = 16'b1010100111011101;
        227: y = 16'b1010100001000001;
        228: y = 16'b1010011010101010;
        229: y = 16'b1010010100011011;
        230: y = 16'b1010001110010010;
        231: y = 16'b1010001000010001;
        232: y = 16'b1010000010010110;
        233: y = 16'b1001111100100011;
        234: y = 16'b1001110110110111;
        235: y = 16'b1001110001010010;
        236: y = 16'b1001101011110101;
        237: y = 16'b1001100110100000;
        238: y = 16'b1001100001010010;
        239: y = 16'b1001011100001100;
        240: y = 16'b1001010111001110;
        241: y = 16'b1001010010011000;
        242: y = 16'b1001001101101010;
        243: y = 16'b1001001001000100;
        244: y = 16'b1001000100100111;
        245: y = 16'b1001000000010010;
        246: y = 16'b1000111100000101;
        247: y = 16'b1000111000000001;
        248: y = 16'b1000110100000110;
        249: y = 16'b1000110000010011;
        250: y = 16'b1000101100101001;
        251: y = 16'b1000101001001000;
        252: y = 16'b1000100101101111;
        253: y = 16'b1000100010100000;
        254: y = 16'b1000011111011001;
        255: y = 16'b1000011100011100;
        256: y = 16'b1000011001101000;
        257: y = 16'b1000010110111101;
        258: y = 16'b1000010100011011;
        259: y = 16'b1000010010000010;
        260: y = 16'b1000001111110011;
        261: y = 16'b1000001101101101;
        262: y = 16'b1000001011110001;
        263: y = 16'b1000001001111101;
        264: y = 16'b1000001000010100;
        265: y = 16'b1000000110110100;
        266: y = 16'b1000000101011101;
        267: y = 16'b1000000100010000;
        268: y = 16'b1000000011001101;
        269: y = 16'b1000000010010011;
        270: y = 16'b1000000001100011;
        271: y = 16'b1000000000111100;
        272: y = 16'b1000000000011111;
        273: y = 16'b1000000000001100;
        274: y = 16'b1000000000000010;
        275: y = 16'b1000000000000010;
        276: y = 16'b1000000000001100;
        277: y = 16'b1000000000011111;
        278: y = 16'b1000000000111100;
        279: y = 16'b1000000001100011;
        280: y = 16'b1000000010010011;
        281: y = 16'b1000000011001101;
        282: y = 16'b1000000100010000;
        283: y = 16'b1000000101011101;
        284: y = 16'b1000000110110100;
        285: y = 16'b1000001000010100;
        286: y = 16'b1000001001111101;
        287: y = 16'b1000001011110001;
        288: y = 16'b1000001101101101;
        289: y = 16'b1000001111110011;
        290: y = 16'b1000010010000010;
        291: y = 16'b1000010100011011;
        292: y = 16'b1000010110111101;
        293: y = 16'b1000011001101000;
        294: y = 16'b1000011100011100;
        295: y = 16'b1000011111011001;
        296: y = 16'b1000100010100000;
        297: y = 16'b1000100101101111;
        298: y = 16'b1000101001001000;
        299: y = 16'b1000101100101001;
        300: y = 16'b1000110000010011;
        301: y = 16'b1000110100000110;
        302: y = 16'b1000111000000001;
        303: y = 16'b1000111100000101;
        304: y = 16'b1001000000010010;
        305: y = 16'b1001000100100111;
        306: y = 16'b1001001001000100;
        307: y = 16'b1001001101101010;
        308: y = 16'b1001010010011000;
        309: y = 16'b1001010111001110;
        310: y = 16'b1001011100001100;
        311: y = 16'b1001100001010010;
        312: y = 16'b1001100110100000;
        313: y = 16'b1001101011110101;
        314: y = 16'b1001110001010010;
        315: y = 16'b1001110110110111;
        316: y = 16'b1001111100100011;
        317: y = 16'b1010000010010110;
        318: y = 16'b1010001000010001;
        319: y = 16'b1010001110010010;
        320: y = 16'b1010010100011011;
        321: y = 16'b1010011010101010;
        322: y = 16'b1010100001000001;
        323: y = 16'b1010100111011101;
        324: y = 16'b1010101110000001;
        325: y = 16'b1010110100101010;
        326: y = 16'b1010111011011010;
        327: y = 16'b1011000010010000;
        328: y = 16'b1011001001001101;
        329: y = 16'b1011010000001110;
        330: y = 16'b1011010111010110;
        331: y = 16'b1011011110100011;
        332: y = 16'b1011100101110110;
        333: y = 16'b1011101101001110;
        334: y = 16'b1011110100101011;
        335: y = 16'b1011111100001110;
        336: y = 16'b1100000011110101;
        337: y = 16'b1100001011100001;
        338: y = 16'b1100010011010001;
        339: y = 16'b1100011011000110;
        340: y = 16'b1100100010111111;
        341: y = 16'b1100101010111101;
        342: y = 16'b1100110010111110;
        343: y = 16'b1100111011000100;
        344: y = 16'b1101000011001101;
        345: y = 16'b1101001011011001;
        346: y = 16'b1101010011101001;
        347: y = 16'b1101011011111101;
        348: y = 16'b1101100100010011;
        349: y = 16'b1101101100101100;
        350: y = 16'b1101110101001000;
        351: y = 16'b1101111101100111;
        352: y = 16'b1110000110001000;
        353: y = 16'b1110001110101100;
        354: y = 16'b1110010111010001;
        355: y = 16'b1110011111111001;
        356: y = 16'b1110101000100010;
        357: y = 16'b1110110001001101;
        358: y = 16'b1110111001111010;
        359: y = 16'b1111000010101000;
        360: y = 16'b1111001011010111;
        361: y = 16'b1111010100000111;
        362: y = 16'b1111011100111000;
        363: y = 16'b1111100101101001;
        364: y = 16'b1111101110011011;
        365: y = 16'b1111110111001110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=277.18Hz, Fs=96000Hz, 16-bit

module lut_Cs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 345;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001001010011;
        2: y = 16'b0000010010100110;
        3: y = 16'b0000011011111000;
        4: y = 16'b0000100101001010;
        5: y = 16'b0000101110011011;
        6: y = 16'b0000110111101011;
        7: y = 16'b0001000000111010;
        8: y = 16'b0001001010001000;
        9: y = 16'b0001010011010011;
        10: y = 16'b0001011100011110;
        11: y = 16'b0001100101100110;
        12: y = 16'b0001101110101100;
        13: y = 16'b0001110111110000;
        14: y = 16'b0010000000110001;
        15: y = 16'b0010001001110000;
        16: y = 16'b0010010010101011;
        17: y = 16'b0010011011100100;
        18: y = 16'b0010100100011001;
        19: y = 16'b0010101101001011;
        20: y = 16'b0010110101111001;
        21: y = 16'b0010111110100011;
        22: y = 16'b0011000111001001;
        23: y = 16'b0011001111101011;
        24: y = 16'b0011011000001001;
        25: y = 16'b0011100000100010;
        26: y = 16'b0011101000110110;
        27: y = 16'b0011110001000110;
        28: y = 16'b0011111001010000;
        29: y = 16'b0100000001010101;
        30: y = 16'b0100001001010101;
        31: y = 16'b0100010001001111;
        32: y = 16'b0100011001000011;
        33: y = 16'b0100100000110010;
        34: y = 16'b0100101000011010;
        35: y = 16'b0100101111111100;
        36: y = 16'b0100110111011000;
        37: y = 16'b0100111110101101;
        38: y = 16'b0101000101111011;
        39: y = 16'b0101001101000010;
        40: y = 16'b0101010100000011;
        41: y = 16'b0101011010111100;
        42: y = 16'b0101100001101110;
        43: y = 16'b0101101000011000;
        44: y = 16'b0101101110111011;
        45: y = 16'b0101110101010110;
        46: y = 16'b0101111011101001;
        47: y = 16'b0110000001110101;
        48: y = 16'b0110000111111000;
        49: y = 16'b0110001101110010;
        50: y = 16'b0110010011100101;
        51: y = 16'b0110011001001111;
        52: y = 16'b0110011110110000;
        53: y = 16'b0110100100001000;
        54: y = 16'b0110101001011000;
        55: y = 16'b0110101110011111;
        56: y = 16'b0110110011011100;
        57: y = 16'b0110111000010001;
        58: y = 16'b0110111100111100;
        59: y = 16'b0111000001011101;
        60: y = 16'b0111000101110110;
        61: y = 16'b0111001010000100;
        62: y = 16'b0111001110001001;
        63: y = 16'b0111010010000100;
        64: y = 16'b0111010101110110;
        65: y = 16'b0111011001011101;
        66: y = 16'b0111011100111011;
        67: y = 16'b0111100000001110;
        68: y = 16'b0111100011010111;
        69: y = 16'b0111100110010110;
        70: y = 16'b0111101001001011;
        71: y = 16'b0111101011110110;
        72: y = 16'b0111101110010110;
        73: y = 16'b0111110000101011;
        74: y = 16'b0111110010110110;
        75: y = 16'b0111110100110111;
        76: y = 16'b0111110110101101;
        77: y = 16'b0111111000011001;
        78: y = 16'b0111111001111001;
        79: y = 16'b0111111011010000;
        80: y = 16'b0111111100011011;
        81: y = 16'b0111111101011100;
        82: y = 16'b0111111110010010;
        83: y = 16'b0111111110111101;
        84: y = 16'b0111111111011101;
        85: y = 16'b0111111111110011;
        86: y = 16'b0111111111111110;
        87: y = 16'b0111111111111110;
        88: y = 16'b0111111111110011;
        89: y = 16'b0111111111011101;
        90: y = 16'b0111111110111101;
        91: y = 16'b0111111110010010;
        92: y = 16'b0111111101011100;
        93: y = 16'b0111111100011011;
        94: y = 16'b0111111011010000;
        95: y = 16'b0111111001111001;
        96: y = 16'b0111111000011001;
        97: y = 16'b0111110110101101;
        98: y = 16'b0111110100110111;
        99: y = 16'b0111110010110110;
        100: y = 16'b0111110000101011;
        101: y = 16'b0111101110010110;
        102: y = 16'b0111101011110110;
        103: y = 16'b0111101001001011;
        104: y = 16'b0111100110010110;
        105: y = 16'b0111100011010111;
        106: y = 16'b0111100000001110;
        107: y = 16'b0111011100111011;
        108: y = 16'b0111011001011101;
        109: y = 16'b0111010101110110;
        110: y = 16'b0111010010000100;
        111: y = 16'b0111001110001001;
        112: y = 16'b0111001010000100;
        113: y = 16'b0111000101110110;
        114: y = 16'b0111000001011101;
        115: y = 16'b0110111100111100;
        116: y = 16'b0110111000010001;
        117: y = 16'b0110110011011100;
        118: y = 16'b0110101110011111;
        119: y = 16'b0110101001011000;
        120: y = 16'b0110100100001000;
        121: y = 16'b0110011110110000;
        122: y = 16'b0110011001001111;
        123: y = 16'b0110010011100101;
        124: y = 16'b0110001101110010;
        125: y = 16'b0110000111111000;
        126: y = 16'b0110000001110101;
        127: y = 16'b0101111011101001;
        128: y = 16'b0101110101010110;
        129: y = 16'b0101101110111011;
        130: y = 16'b0101101000011000;
        131: y = 16'b0101100001101110;
        132: y = 16'b0101011010111100;
        133: y = 16'b0101010100000011;
        134: y = 16'b0101001101000010;
        135: y = 16'b0101000101111011;
        136: y = 16'b0100111110101101;
        137: y = 16'b0100110111011000;
        138: y = 16'b0100101111111100;
        139: y = 16'b0100101000011010;
        140: y = 16'b0100100000110010;
        141: y = 16'b0100011001000011;
        142: y = 16'b0100010001001111;
        143: y = 16'b0100001001010101;
        144: y = 16'b0100000001010101;
        145: y = 16'b0011111001010000;
        146: y = 16'b0011110001000110;
        147: y = 16'b0011101000110110;
        148: y = 16'b0011100000100010;
        149: y = 16'b0011011000001001;
        150: y = 16'b0011001111101011;
        151: y = 16'b0011000111001001;
        152: y = 16'b0010111110100011;
        153: y = 16'b0010110101111001;
        154: y = 16'b0010101101001011;
        155: y = 16'b0010100100011001;
        156: y = 16'b0010011011100100;
        157: y = 16'b0010010010101011;
        158: y = 16'b0010001001110000;
        159: y = 16'b0010000000110001;
        160: y = 16'b0001110111110000;
        161: y = 16'b0001101110101100;
        162: y = 16'b0001100101100110;
        163: y = 16'b0001011100011110;
        164: y = 16'b0001010011010011;
        165: y = 16'b0001001010001000;
        166: y = 16'b0001000000111010;
        167: y = 16'b0000110111101011;
        168: y = 16'b0000101110011011;
        169: y = 16'b0000100101001010;
        170: y = 16'b0000011011111000;
        171: y = 16'b0000010010100110;
        172: y = 16'b0000001001010011;
        173: y = 16'b0000000000000000;
        174: y = 16'b1111110110101101;
        175: y = 16'b1111101101011010;
        176: y = 16'b1111100100001000;
        177: y = 16'b1111011010110110;
        178: y = 16'b1111010001100101;
        179: y = 16'b1111001000010101;
        180: y = 16'b1110111111000110;
        181: y = 16'b1110110101111000;
        182: y = 16'b1110101100101101;
        183: y = 16'b1110100011100010;
        184: y = 16'b1110011010011010;
        185: y = 16'b1110010001010100;
        186: y = 16'b1110001000010000;
        187: y = 16'b1101111111001111;
        188: y = 16'b1101110110010000;
        189: y = 16'b1101101101010101;
        190: y = 16'b1101100100011100;
        191: y = 16'b1101011011100111;
        192: y = 16'b1101010010110101;
        193: y = 16'b1101001010000111;
        194: y = 16'b1101000001011101;
        195: y = 16'b1100111000110111;
        196: y = 16'b1100110000010101;
        197: y = 16'b1100100111110111;
        198: y = 16'b1100011111011110;
        199: y = 16'b1100010111001010;
        200: y = 16'b1100001110111010;
        201: y = 16'b1100000110110000;
        202: y = 16'b1011111110101011;
        203: y = 16'b1011110110101011;
        204: y = 16'b1011101110110001;
        205: y = 16'b1011100110111101;
        206: y = 16'b1011011111001110;
        207: y = 16'b1011010111100110;
        208: y = 16'b1011010000000100;
        209: y = 16'b1011001000101000;
        210: y = 16'b1011000001010011;
        211: y = 16'b1010111010000101;
        212: y = 16'b1010110010111110;
        213: y = 16'b1010101011111101;
        214: y = 16'b1010100101000100;
        215: y = 16'b1010011110010010;
        216: y = 16'b1010010111101000;
        217: y = 16'b1010010001000101;
        218: y = 16'b1010001010101010;
        219: y = 16'b1010000100010111;
        220: y = 16'b1001111110001011;
        221: y = 16'b1001111000001000;
        222: y = 16'b1001110010001110;
        223: y = 16'b1001101100011011;
        224: y = 16'b1001100110110001;
        225: y = 16'b1001100001010000;
        226: y = 16'b1001011011111000;
        227: y = 16'b1001010110101000;
        228: y = 16'b1001010001100001;
        229: y = 16'b1001001100100100;
        230: y = 16'b1001000111101111;
        231: y = 16'b1001000011000100;
        232: y = 16'b1000111110100011;
        233: y = 16'b1000111010001010;
        234: y = 16'b1000110101111100;
        235: y = 16'b1000110001110111;
        236: y = 16'b1000101101111100;
        237: y = 16'b1000101010001010;
        238: y = 16'b1000100110100011;
        239: y = 16'b1000100011000101;
        240: y = 16'b1000011111110010;
        241: y = 16'b1000011100101001;
        242: y = 16'b1000011001101010;
        243: y = 16'b1000010110110101;
        244: y = 16'b1000010100001010;
        245: y = 16'b1000010001101010;
        246: y = 16'b1000001111010101;
        247: y = 16'b1000001101001010;
        248: y = 16'b1000001011001001;
        249: y = 16'b1000001001010011;
        250: y = 16'b1000000111100111;
        251: y = 16'b1000000110000111;
        252: y = 16'b1000000100110000;
        253: y = 16'b1000000011100101;
        254: y = 16'b1000000010100100;
        255: y = 16'b1000000001101110;
        256: y = 16'b1000000001000011;
        257: y = 16'b1000000000100011;
        258: y = 16'b1000000000001101;
        259: y = 16'b1000000000000010;
        260: y = 16'b1000000000000010;
        261: y = 16'b1000000000001101;
        262: y = 16'b1000000000100011;
        263: y = 16'b1000000001000011;
        264: y = 16'b1000000001101110;
        265: y = 16'b1000000010100100;
        266: y = 16'b1000000011100101;
        267: y = 16'b1000000100110000;
        268: y = 16'b1000000110000111;
        269: y = 16'b1000000111100111;
        270: y = 16'b1000001001010011;
        271: y = 16'b1000001011001001;
        272: y = 16'b1000001101001010;
        273: y = 16'b1000001111010101;
        274: y = 16'b1000010001101010;
        275: y = 16'b1000010100001010;
        276: y = 16'b1000010110110101;
        277: y = 16'b1000011001101010;
        278: y = 16'b1000011100101001;
        279: y = 16'b1000011111110010;
        280: y = 16'b1000100011000101;
        281: y = 16'b1000100110100011;
        282: y = 16'b1000101010001010;
        283: y = 16'b1000101101111100;
        284: y = 16'b1000110001110111;
        285: y = 16'b1000110101111100;
        286: y = 16'b1000111010001010;
        287: y = 16'b1000111110100011;
        288: y = 16'b1001000011000100;
        289: y = 16'b1001000111101111;
        290: y = 16'b1001001100100100;
        291: y = 16'b1001010001100001;
        292: y = 16'b1001010110101000;
        293: y = 16'b1001011011111000;
        294: y = 16'b1001100001010000;
        295: y = 16'b1001100110110001;
        296: y = 16'b1001101100011011;
        297: y = 16'b1001110010001110;
        298: y = 16'b1001111000001000;
        299: y = 16'b1001111110001011;
        300: y = 16'b1010000100010111;
        301: y = 16'b1010001010101010;
        302: y = 16'b1010010001000101;
        303: y = 16'b1010010111101000;
        304: y = 16'b1010011110010010;
        305: y = 16'b1010100101000100;
        306: y = 16'b1010101011111101;
        307: y = 16'b1010110010111110;
        308: y = 16'b1010111010000101;
        309: y = 16'b1011000001010011;
        310: y = 16'b1011001000101000;
        311: y = 16'b1011010000000100;
        312: y = 16'b1011010111100110;
        313: y = 16'b1011011111001110;
        314: y = 16'b1011100110111101;
        315: y = 16'b1011101110110001;
        316: y = 16'b1011110110101011;
        317: y = 16'b1011111110101011;
        318: y = 16'b1100000110110000;
        319: y = 16'b1100001110111010;
        320: y = 16'b1100010111001010;
        321: y = 16'b1100011111011110;
        322: y = 16'b1100100111110111;
        323: y = 16'b1100110000010101;
        324: y = 16'b1100111000110111;
        325: y = 16'b1101000001011101;
        326: y = 16'b1101001010000111;
        327: y = 16'b1101010010110101;
        328: y = 16'b1101011011100111;
        329: y = 16'b1101100100011100;
        330: y = 16'b1101101101010101;
        331: y = 16'b1101110110010000;
        332: y = 16'b1101111111001111;
        333: y = 16'b1110001000010000;
        334: y = 16'b1110010001010100;
        335: y = 16'b1110011010011010;
        336: y = 16'b1110100011100010;
        337: y = 16'b1110101100101101;
        338: y = 16'b1110110101111000;
        339: y = 16'b1110111111000110;
        340: y = 16'b1111001000010101;
        341: y = 16'b1111010001100101;
        342: y = 16'b1111011010110110;
        343: y = 16'b1111100100001000;
        344: y = 16'b1111101101011010;
        345: y = 16'b1111110110101101;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=293.66Hz, Fs=96000Hz, 16-bit

module lut_D
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 325;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001001110111;
        2: y = 16'b0000010011101111;
        3: y = 16'b0000011101100110;
        4: y = 16'b0000100111011100;
        5: y = 16'b0000110001010001;
        6: y = 16'b0000111011000101;
        7: y = 16'b0001000100110111;
        8: y = 16'b0001001110101000;
        9: y = 16'b0001011000010111;
        10: y = 16'b0001100010000100;
        11: y = 16'b0001101011101111;
        12: y = 16'b0001110101010111;
        13: y = 16'b0001111110111100;
        14: y = 16'b0010001000011111;
        15: y = 16'b0010010001111110;
        16: y = 16'b0010011011011001;
        17: y = 16'b0010100100110001;
        18: y = 16'b0010101110000101;
        19: y = 16'b0010110111010101;
        20: y = 16'b0011000000100000;
        21: y = 16'b0011001001100111;
        22: y = 16'b0011010010101001;
        23: y = 16'b0011011011100110;
        24: y = 16'b0011100100011110;
        25: y = 16'b0011101101010001;
        26: y = 16'b0011110101111101;
        27: y = 16'b0011111110100100;
        28: y = 16'b0100000111000101;
        29: y = 16'b0100001111100000;
        30: y = 16'b0100010111110100;
        31: y = 16'b0100100000000001;
        32: y = 16'b0100101000001000;
        33: y = 16'b0100110000001000;
        34: y = 16'b0100111000000000;
        35: y = 16'b0100111111110001;
        36: y = 16'b0101000111011011;
        37: y = 16'b0101001110111100;
        38: y = 16'b0101010110010110;
        39: y = 16'b0101011101100111;
        40: y = 16'b0101100100110000;
        41: y = 16'b0101101011110001;
        42: y = 16'b0101110010101001;
        43: y = 16'b0101111001011000;
        44: y = 16'b0101111111111111;
        45: y = 16'b0110000110011100;
        46: y = 16'b0110001100110000;
        47: y = 16'b0110010010111010;
        48: y = 16'b0110011000111011;
        49: y = 16'b0110011110110010;
        50: y = 16'b0110100100011111;
        51: y = 16'b0110101010000011;
        52: y = 16'b0110101111011100;
        53: y = 16'b0110110100101011;
        54: y = 16'b0110111001101111;
        55: y = 16'b0110111110101001;
        56: y = 16'b0111000011011001;
        57: y = 16'b0111000111111101;
        58: y = 16'b0111001100010111;
        59: y = 16'b0111010000100110;
        60: y = 16'b0111010100101010;
        61: y = 16'b0111011000100010;
        62: y = 16'b0111011100010000;
        63: y = 16'b0111011111110010;
        64: y = 16'b0111100011001001;
        65: y = 16'b0111100110010100;
        66: y = 16'b0111101001010100;
        67: y = 16'b0111101100001000;
        68: y = 16'b0111101110110000;
        69: y = 16'b0111110001001101;
        70: y = 16'b0111110011011101;
        71: y = 16'b0111110101100010;
        72: y = 16'b0111110111011011;
        73: y = 16'b0111111001001000;
        74: y = 16'b0111111010101001;
        75: y = 16'b0111111011111110;
        76: y = 16'b0111111101000111;
        77: y = 16'b0111111110000100;
        78: y = 16'b0111111110110100;
        79: y = 16'b0111111111011001;
        80: y = 16'b0111111111110001;
        81: y = 16'b0111111111111101;
        82: y = 16'b0111111111111101;
        83: y = 16'b0111111111110001;
        84: y = 16'b0111111111011001;
        85: y = 16'b0111111110110100;
        86: y = 16'b0111111110000100;
        87: y = 16'b0111111101000111;
        88: y = 16'b0111111011111110;
        89: y = 16'b0111111010101001;
        90: y = 16'b0111111001001000;
        91: y = 16'b0111110111011011;
        92: y = 16'b0111110101100010;
        93: y = 16'b0111110011011101;
        94: y = 16'b0111110001001101;
        95: y = 16'b0111101110110000;
        96: y = 16'b0111101100001000;
        97: y = 16'b0111101001010100;
        98: y = 16'b0111100110010100;
        99: y = 16'b0111100011001001;
        100: y = 16'b0111011111110010;
        101: y = 16'b0111011100010000;
        102: y = 16'b0111011000100010;
        103: y = 16'b0111010100101010;
        104: y = 16'b0111010000100110;
        105: y = 16'b0111001100010111;
        106: y = 16'b0111000111111101;
        107: y = 16'b0111000011011001;
        108: y = 16'b0110111110101001;
        109: y = 16'b0110111001101111;
        110: y = 16'b0110110100101011;
        111: y = 16'b0110101111011100;
        112: y = 16'b0110101010000011;
        113: y = 16'b0110100100011111;
        114: y = 16'b0110011110110010;
        115: y = 16'b0110011000111011;
        116: y = 16'b0110010010111010;
        117: y = 16'b0110001100110000;
        118: y = 16'b0110000110011100;
        119: y = 16'b0101111111111111;
        120: y = 16'b0101111001011000;
        121: y = 16'b0101110010101001;
        122: y = 16'b0101101011110001;
        123: y = 16'b0101100100110000;
        124: y = 16'b0101011101100111;
        125: y = 16'b0101010110010110;
        126: y = 16'b0101001110111100;
        127: y = 16'b0101000111011011;
        128: y = 16'b0100111111110001;
        129: y = 16'b0100111000000000;
        130: y = 16'b0100110000001000;
        131: y = 16'b0100101000001000;
        132: y = 16'b0100100000000001;
        133: y = 16'b0100010111110100;
        134: y = 16'b0100001111100000;
        135: y = 16'b0100000111000101;
        136: y = 16'b0011111110100100;
        137: y = 16'b0011110101111101;
        138: y = 16'b0011101101010001;
        139: y = 16'b0011100100011110;
        140: y = 16'b0011011011100110;
        141: y = 16'b0011010010101001;
        142: y = 16'b0011001001100111;
        143: y = 16'b0011000000100000;
        144: y = 16'b0010110111010101;
        145: y = 16'b0010101110000101;
        146: y = 16'b0010100100110001;
        147: y = 16'b0010011011011001;
        148: y = 16'b0010010001111110;
        149: y = 16'b0010001000011111;
        150: y = 16'b0001111110111100;
        151: y = 16'b0001110101010111;
        152: y = 16'b0001101011101111;
        153: y = 16'b0001100010000100;
        154: y = 16'b0001011000010111;
        155: y = 16'b0001001110101000;
        156: y = 16'b0001000100110111;
        157: y = 16'b0000111011000101;
        158: y = 16'b0000110001010001;
        159: y = 16'b0000100111011100;
        160: y = 16'b0000011101100110;
        161: y = 16'b0000010011101111;
        162: y = 16'b0000001001110111;
        163: y = 16'b0000000000000000;
        164: y = 16'b1111110110001001;
        165: y = 16'b1111101100010001;
        166: y = 16'b1111100010011010;
        167: y = 16'b1111011000100100;
        168: y = 16'b1111001110101111;
        169: y = 16'b1111000100111011;
        170: y = 16'b1110111011001001;
        171: y = 16'b1110110001011000;
        172: y = 16'b1110100111101001;
        173: y = 16'b1110011101111100;
        174: y = 16'b1110010100010001;
        175: y = 16'b1110001010101001;
        176: y = 16'b1110000001000100;
        177: y = 16'b1101110111100001;
        178: y = 16'b1101101110000010;
        179: y = 16'b1101100100100111;
        180: y = 16'b1101011011001111;
        181: y = 16'b1101010001111011;
        182: y = 16'b1101001000101011;
        183: y = 16'b1100111111100000;
        184: y = 16'b1100110110011001;
        185: y = 16'b1100101101010111;
        186: y = 16'b1100100100011010;
        187: y = 16'b1100011011100010;
        188: y = 16'b1100010010101111;
        189: y = 16'b1100001010000011;
        190: y = 16'b1100000001011100;
        191: y = 16'b1011111000111011;
        192: y = 16'b1011110000100000;
        193: y = 16'b1011101000001100;
        194: y = 16'b1011011111111111;
        195: y = 16'b1011010111111000;
        196: y = 16'b1011001111111000;
        197: y = 16'b1011001000000000;
        198: y = 16'b1011000000001111;
        199: y = 16'b1010111000100101;
        200: y = 16'b1010110001000100;
        201: y = 16'b1010101001101010;
        202: y = 16'b1010100010011001;
        203: y = 16'b1010011011010000;
        204: y = 16'b1010010100001111;
        205: y = 16'b1010001101010111;
        206: y = 16'b1010000110101000;
        207: y = 16'b1010000000000001;
        208: y = 16'b1001111001100100;
        209: y = 16'b1001110011010000;
        210: y = 16'b1001101101000110;
        211: y = 16'b1001100111000101;
        212: y = 16'b1001100001001110;
        213: y = 16'b1001011011100001;
        214: y = 16'b1001010101111101;
        215: y = 16'b1001010000100100;
        216: y = 16'b1001001011010101;
        217: y = 16'b1001000110010001;
        218: y = 16'b1001000001010111;
        219: y = 16'b1000111100100111;
        220: y = 16'b1000111000000011;
        221: y = 16'b1000110011101001;
        222: y = 16'b1000101111011010;
        223: y = 16'b1000101011010110;
        224: y = 16'b1000100111011110;
        225: y = 16'b1000100011110000;
        226: y = 16'b1000100000001110;
        227: y = 16'b1000011100110111;
        228: y = 16'b1000011001101100;
        229: y = 16'b1000010110101100;
        230: y = 16'b1000010011111000;
        231: y = 16'b1000010001010000;
        232: y = 16'b1000001110110011;
        233: y = 16'b1000001100100011;
        234: y = 16'b1000001010011110;
        235: y = 16'b1000001000100101;
        236: y = 16'b1000000110111000;
        237: y = 16'b1000000101010111;
        238: y = 16'b1000000100000010;
        239: y = 16'b1000000010111001;
        240: y = 16'b1000000001111100;
        241: y = 16'b1000000001001100;
        242: y = 16'b1000000000100111;
        243: y = 16'b1000000000001111;
        244: y = 16'b1000000000000011;
        245: y = 16'b1000000000000011;
        246: y = 16'b1000000000001111;
        247: y = 16'b1000000000100111;
        248: y = 16'b1000000001001100;
        249: y = 16'b1000000001111100;
        250: y = 16'b1000000010111001;
        251: y = 16'b1000000100000010;
        252: y = 16'b1000000101010111;
        253: y = 16'b1000000110111000;
        254: y = 16'b1000001000100101;
        255: y = 16'b1000001010011110;
        256: y = 16'b1000001100100011;
        257: y = 16'b1000001110110011;
        258: y = 16'b1000010001010000;
        259: y = 16'b1000010011111000;
        260: y = 16'b1000010110101100;
        261: y = 16'b1000011001101100;
        262: y = 16'b1000011100110111;
        263: y = 16'b1000100000001110;
        264: y = 16'b1000100011110000;
        265: y = 16'b1000100111011110;
        266: y = 16'b1000101011010110;
        267: y = 16'b1000101111011010;
        268: y = 16'b1000110011101001;
        269: y = 16'b1000111000000011;
        270: y = 16'b1000111100100111;
        271: y = 16'b1001000001010111;
        272: y = 16'b1001000110010001;
        273: y = 16'b1001001011010101;
        274: y = 16'b1001010000100100;
        275: y = 16'b1001010101111101;
        276: y = 16'b1001011011100001;
        277: y = 16'b1001100001001110;
        278: y = 16'b1001100111000101;
        279: y = 16'b1001101101000110;
        280: y = 16'b1001110011010000;
        281: y = 16'b1001111001100100;
        282: y = 16'b1010000000000001;
        283: y = 16'b1010000110101000;
        284: y = 16'b1010001101010111;
        285: y = 16'b1010010100001111;
        286: y = 16'b1010011011010000;
        287: y = 16'b1010100010011001;
        288: y = 16'b1010101001101010;
        289: y = 16'b1010110001000100;
        290: y = 16'b1010111000100101;
        291: y = 16'b1011000000001111;
        292: y = 16'b1011001000000000;
        293: y = 16'b1011001111111000;
        294: y = 16'b1011010111111000;
        295: y = 16'b1011011111111111;
        296: y = 16'b1011101000001100;
        297: y = 16'b1011110000100000;
        298: y = 16'b1011111000111011;
        299: y = 16'b1100000001011100;
        300: y = 16'b1100001010000011;
        301: y = 16'b1100010010101111;
        302: y = 16'b1100011011100010;
        303: y = 16'b1100100100011010;
        304: y = 16'b1100101101010111;
        305: y = 16'b1100110110011001;
        306: y = 16'b1100111111100000;
        307: y = 16'b1101001000101011;
        308: y = 16'b1101010001111011;
        309: y = 16'b1101011011001111;
        310: y = 16'b1101100100100111;
        311: y = 16'b1101101110000010;
        312: y = 16'b1101110111100001;
        313: y = 16'b1110000001000100;
        314: y = 16'b1110001010101001;
        315: y = 16'b1110010100010001;
        316: y = 16'b1110011101111100;
        317: y = 16'b1110100111101001;
        318: y = 16'b1110110001011000;
        319: y = 16'b1110111011001001;
        320: y = 16'b1111000100111011;
        321: y = 16'b1111001110101111;
        322: y = 16'b1111011000100100;
        323: y = 16'b1111100010011010;
        324: y = 16'b1111101100010001;
        325: y = 16'b1111110110001001;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=311.13Hz, Fs=96000Hz, 16-bit

module lut_Ds
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 307;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001010011100;
        2: y = 16'b0000010100111001;
        3: y = 16'b0000011111010100;
        4: y = 16'b0000101001101111;
        5: y = 16'b0000110100001000;
        6: y = 16'b0000111110100001;
        7: y = 16'b0001001000110111;
        8: y = 16'b0001010011001100;
        9: y = 16'b0001011101011110;
        10: y = 16'b0001100111101110;
        11: y = 16'b0001110001111011;
        12: y = 16'b0001111100000101;
        13: y = 16'b0010000110001100;
        14: y = 16'b0010010000010000;
        15: y = 16'b0010011010001111;
        16: y = 16'b0010100100001010;
        17: y = 16'b0010101110000001;
        18: y = 16'b0010110111110011;
        19: y = 16'b0011000001100001;
        20: y = 16'b0011001011001001;
        21: y = 16'b0011010100101100;
        22: y = 16'b0011011110001001;
        23: y = 16'b0011100111100000;
        24: y = 16'b0011110000110001;
        25: y = 16'b0011111001111100;
        26: y = 16'b0100000011000000;
        27: y = 16'b0100001011111101;
        28: y = 16'b0100010100110011;
        29: y = 16'b0100011101100010;
        30: y = 16'b0100100110001001;
        31: y = 16'b0100101110101000;
        32: y = 16'b0100110110111111;
        33: y = 16'b0100111111001110;
        34: y = 16'b0101000111010100;
        35: y = 16'b0101001111010010;
        36: y = 16'b0101010111000110;
        37: y = 16'b0101011110110010;
        38: y = 16'b0101100110010100;
        39: y = 16'b0101101101101101;
        40: y = 16'b0101110100111100;
        41: y = 16'b0101111100000001;
        42: y = 16'b0110000010111100;
        43: y = 16'b0110001001101100;
        44: y = 16'b0110010000010010;
        45: y = 16'b0110010110101110;
        46: y = 16'b0110011100111110;
        47: y = 16'b0110100011000100;
        48: y = 16'b0110101000111110;
        49: y = 16'b0110101110101101;
        50: y = 16'b0110110100010001;
        51: y = 16'b0110111001101001;
        52: y = 16'b0110111110110101;
        53: y = 16'b0111000011110110;
        54: y = 16'b0111001000101010;
        55: y = 16'b0111001101010010;
        56: y = 16'b0111010001101110;
        57: y = 16'b0111010101111101;
        58: y = 16'b0111011010000000;
        59: y = 16'b0111011101110111;
        60: y = 16'b0111100001100000;
        61: y = 16'b0111100100111101;
        62: y = 16'b0111101000001101;
        63: y = 16'b0111101011010000;
        64: y = 16'b0111101110000101;
        65: y = 16'b0111110000101110;
        66: y = 16'b0111110011001001;
        67: y = 16'b0111110101011000;
        68: y = 16'b0111110111011000;
        69: y = 16'b0111111001001100;
        70: y = 16'b0111111010110001;
        71: y = 16'b0111111100001010;
        72: y = 16'b0111111101010101;
        73: y = 16'b0111111110010010;
        74: y = 16'b0111111111000010;
        75: y = 16'b0111111111100100;
        76: y = 16'b0111111111111000;
        77: y = 16'b0111111111111111;
        78: y = 16'b0111111111111000;
        79: y = 16'b0111111111100100;
        80: y = 16'b0111111111000010;
        81: y = 16'b0111111110010010;
        82: y = 16'b0111111101010101;
        83: y = 16'b0111111100001010;
        84: y = 16'b0111111010110001;
        85: y = 16'b0111111001001100;
        86: y = 16'b0111110111011000;
        87: y = 16'b0111110101011000;
        88: y = 16'b0111110011001001;
        89: y = 16'b0111110000101110;
        90: y = 16'b0111101110000101;
        91: y = 16'b0111101011010000;
        92: y = 16'b0111101000001101;
        93: y = 16'b0111100100111101;
        94: y = 16'b0111100001100000;
        95: y = 16'b0111011101110111;
        96: y = 16'b0111011010000000;
        97: y = 16'b0111010101111101;
        98: y = 16'b0111010001101110;
        99: y = 16'b0111001101010010;
        100: y = 16'b0111001000101010;
        101: y = 16'b0111000011110110;
        102: y = 16'b0110111110110101;
        103: y = 16'b0110111001101001;
        104: y = 16'b0110110100010001;
        105: y = 16'b0110101110101101;
        106: y = 16'b0110101000111110;
        107: y = 16'b0110100011000100;
        108: y = 16'b0110011100111110;
        109: y = 16'b0110010110101110;
        110: y = 16'b0110010000010010;
        111: y = 16'b0110001001101100;
        112: y = 16'b0110000010111100;
        113: y = 16'b0101111100000001;
        114: y = 16'b0101110100111100;
        115: y = 16'b0101101101101101;
        116: y = 16'b0101100110010100;
        117: y = 16'b0101011110110010;
        118: y = 16'b0101010111000110;
        119: y = 16'b0101001111010010;
        120: y = 16'b0101000111010100;
        121: y = 16'b0100111111001110;
        122: y = 16'b0100110110111111;
        123: y = 16'b0100101110101000;
        124: y = 16'b0100100110001001;
        125: y = 16'b0100011101100010;
        126: y = 16'b0100010100110011;
        127: y = 16'b0100001011111101;
        128: y = 16'b0100000011000000;
        129: y = 16'b0011111001111100;
        130: y = 16'b0011110000110001;
        131: y = 16'b0011100111100000;
        132: y = 16'b0011011110001001;
        133: y = 16'b0011010100101100;
        134: y = 16'b0011001011001001;
        135: y = 16'b0011000001100001;
        136: y = 16'b0010110111110011;
        137: y = 16'b0010101110000001;
        138: y = 16'b0010100100001010;
        139: y = 16'b0010011010001111;
        140: y = 16'b0010010000010000;
        141: y = 16'b0010000110001100;
        142: y = 16'b0001111100000101;
        143: y = 16'b0001110001111011;
        144: y = 16'b0001100111101110;
        145: y = 16'b0001011101011110;
        146: y = 16'b0001010011001100;
        147: y = 16'b0001001000110111;
        148: y = 16'b0000111110100001;
        149: y = 16'b0000110100001000;
        150: y = 16'b0000101001101111;
        151: y = 16'b0000011111010100;
        152: y = 16'b0000010100111001;
        153: y = 16'b0000001010011100;
        154: y = 16'b0000000000000000;
        155: y = 16'b1111110101100100;
        156: y = 16'b1111101011000111;
        157: y = 16'b1111100000101100;
        158: y = 16'b1111010110010001;
        159: y = 16'b1111001011111000;
        160: y = 16'b1111000001011111;
        161: y = 16'b1110110111001001;
        162: y = 16'b1110101100110100;
        163: y = 16'b1110100010100010;
        164: y = 16'b1110011000010010;
        165: y = 16'b1110001110000101;
        166: y = 16'b1110000011111011;
        167: y = 16'b1101111001110100;
        168: y = 16'b1101101111110000;
        169: y = 16'b1101100101110001;
        170: y = 16'b1101011011110110;
        171: y = 16'b1101010001111111;
        172: y = 16'b1101001000001101;
        173: y = 16'b1100111110011111;
        174: y = 16'b1100110100110111;
        175: y = 16'b1100101011010100;
        176: y = 16'b1100100001110111;
        177: y = 16'b1100011000100000;
        178: y = 16'b1100001111001111;
        179: y = 16'b1100000110000100;
        180: y = 16'b1011111101000000;
        181: y = 16'b1011110100000011;
        182: y = 16'b1011101011001101;
        183: y = 16'b1011100010011110;
        184: y = 16'b1011011001110111;
        185: y = 16'b1011010001011000;
        186: y = 16'b1011001001000001;
        187: y = 16'b1011000000110010;
        188: y = 16'b1010111000101100;
        189: y = 16'b1010110000101110;
        190: y = 16'b1010101000111010;
        191: y = 16'b1010100001001110;
        192: y = 16'b1010011001101100;
        193: y = 16'b1010010010010011;
        194: y = 16'b1010001011000100;
        195: y = 16'b1010000011111111;
        196: y = 16'b1001111101000100;
        197: y = 16'b1001110110010100;
        198: y = 16'b1001101111101110;
        199: y = 16'b1001101001010010;
        200: y = 16'b1001100011000010;
        201: y = 16'b1001011100111100;
        202: y = 16'b1001010111000010;
        203: y = 16'b1001010001010011;
        204: y = 16'b1001001011101111;
        205: y = 16'b1001000110010111;
        206: y = 16'b1001000001001011;
        207: y = 16'b1000111100001010;
        208: y = 16'b1000110111010110;
        209: y = 16'b1000110010101110;
        210: y = 16'b1000101110010010;
        211: y = 16'b1000101010000011;
        212: y = 16'b1000100110000000;
        213: y = 16'b1000100010001001;
        214: y = 16'b1000011110100000;
        215: y = 16'b1000011011000011;
        216: y = 16'b1000010111110011;
        217: y = 16'b1000010100110000;
        218: y = 16'b1000010001111011;
        219: y = 16'b1000001111010010;
        220: y = 16'b1000001100110111;
        221: y = 16'b1000001010101000;
        222: y = 16'b1000001000101000;
        223: y = 16'b1000000110110100;
        224: y = 16'b1000000101001111;
        225: y = 16'b1000000011110110;
        226: y = 16'b1000000010101011;
        227: y = 16'b1000000001101110;
        228: y = 16'b1000000000111110;
        229: y = 16'b1000000000011100;
        230: y = 16'b1000000000001000;
        231: y = 16'b1000000000000001;
        232: y = 16'b1000000000001000;
        233: y = 16'b1000000000011100;
        234: y = 16'b1000000000111110;
        235: y = 16'b1000000001101110;
        236: y = 16'b1000000010101011;
        237: y = 16'b1000000011110110;
        238: y = 16'b1000000101001111;
        239: y = 16'b1000000110110100;
        240: y = 16'b1000001000101000;
        241: y = 16'b1000001010101000;
        242: y = 16'b1000001100110111;
        243: y = 16'b1000001111010010;
        244: y = 16'b1000010001111011;
        245: y = 16'b1000010100110000;
        246: y = 16'b1000010111110011;
        247: y = 16'b1000011011000011;
        248: y = 16'b1000011110100000;
        249: y = 16'b1000100010001001;
        250: y = 16'b1000100110000000;
        251: y = 16'b1000101010000011;
        252: y = 16'b1000101110010010;
        253: y = 16'b1000110010101110;
        254: y = 16'b1000110111010110;
        255: y = 16'b1000111100001010;
        256: y = 16'b1001000001001011;
        257: y = 16'b1001000110010111;
        258: y = 16'b1001001011101111;
        259: y = 16'b1001010001010011;
        260: y = 16'b1001010111000010;
        261: y = 16'b1001011100111100;
        262: y = 16'b1001100011000010;
        263: y = 16'b1001101001010010;
        264: y = 16'b1001101111101110;
        265: y = 16'b1001110110010100;
        266: y = 16'b1001111101000100;
        267: y = 16'b1010000011111111;
        268: y = 16'b1010001011000100;
        269: y = 16'b1010010010010011;
        270: y = 16'b1010011001101100;
        271: y = 16'b1010100001001110;
        272: y = 16'b1010101000111010;
        273: y = 16'b1010110000101110;
        274: y = 16'b1010111000101100;
        275: y = 16'b1011000000110010;
        276: y = 16'b1011001001000001;
        277: y = 16'b1011010001011000;
        278: y = 16'b1011011001110111;
        279: y = 16'b1011100010011110;
        280: y = 16'b1011101011001101;
        281: y = 16'b1011110100000011;
        282: y = 16'b1011111101000000;
        283: y = 16'b1100000110000100;
        284: y = 16'b1100001111001111;
        285: y = 16'b1100011000100000;
        286: y = 16'b1100100001110111;
        287: y = 16'b1100101011010100;
        288: y = 16'b1100110100110111;
        289: y = 16'b1100111110011111;
        290: y = 16'b1101001000001101;
        291: y = 16'b1101010001111111;
        292: y = 16'b1101011011110110;
        293: y = 16'b1101100101110001;
        294: y = 16'b1101101111110000;
        295: y = 16'b1101111001110100;
        296: y = 16'b1110000011111011;
        297: y = 16'b1110001110000101;
        298: y = 16'b1110011000010010;
        299: y = 16'b1110100010100010;
        300: y = 16'b1110101100110100;
        301: y = 16'b1110110111001001;
        302: y = 16'b1111000001011111;
        303: y = 16'b1111001011111000;
        304: y = 16'b1111010110010001;
        305: y = 16'b1111100000101100;
        306: y = 16'b1111101011000111;
        307: y = 16'b1111110101100100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=329.63Hz, Fs=96000Hz, 16-bit

module lut_E
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 290;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001011000011;
        2: y = 16'b0000010110000111;
        3: y = 16'b0000100001001001;
        4: y = 16'b0000101100001010;
        5: y = 16'b0000110111001011;
        6: y = 16'b0001000010001001;
        7: y = 16'b0001001101000110;
        8: y = 16'b0001011000000000;
        9: y = 16'b0001100010110111;
        10: y = 16'b0001101101101100;
        11: y = 16'b0001111000011101;
        12: y = 16'b0010000011001011;
        13: y = 16'b0010001101110101;
        14: y = 16'b0010011000011011;
        15: y = 16'b0010100010111100;
        16: y = 16'b0010101101011000;
        17: y = 16'b0010110111101111;
        18: y = 16'b0011000010000001;
        19: y = 16'b0011001100001101;
        20: y = 16'b0011010110010010;
        21: y = 16'b0011100000010010;
        22: y = 16'b0011101010001010;
        23: y = 16'b0011110011111100;
        24: y = 16'b0011111101100110;
        25: y = 16'b0100000111001001;
        26: y = 16'b0100010000100100;
        27: y = 16'b0100011001110111;
        28: y = 16'b0100100011000001;
        29: y = 16'b0100101100000011;
        30: y = 16'b0100110100111011;
        31: y = 16'b0100111101101011;
        32: y = 16'b0101000110010001;
        33: y = 16'b0101001110101101;
        34: y = 16'b0101010111000000;
        35: y = 16'b0101011111001000;
        36: y = 16'b0101100111000101;
        37: y = 16'b0101101110111000;
        38: y = 16'b0101110110100000;
        39: y = 16'b0101111101111101;
        40: y = 16'b0110000101001110;
        41: y = 16'b0110001100010100;
        42: y = 16'b0110010011001110;
        43: y = 16'b0110011001111100;
        44: y = 16'b0110100000011110;
        45: y = 16'b0110100110110011;
        46: y = 16'b0110101100111100;
        47: y = 16'b0110110010111000;
        48: y = 16'b0110111000100111;
        49: y = 16'b0110111110001000;
        50: y = 16'b0111000011011101;
        51: y = 16'b0111001000100100;
        52: y = 16'b0111001101011101;
        53: y = 16'b0111010010001001;
        54: y = 16'b0111010110100110;
        55: y = 16'b0111011010110110;
        56: y = 16'b0111011110110111;
        57: y = 16'b0111100010101010;
        58: y = 16'b0111100110001111;
        59: y = 16'b0111101001100110;
        60: y = 16'b0111101100101101;
        61: y = 16'b0111101111100110;
        62: y = 16'b0111110010010000;
        63: y = 16'b0111110100101100;
        64: y = 16'b0111110110111000;
        65: y = 16'b0111111000110101;
        66: y = 16'b0111111010100100;
        67: y = 16'b0111111100000011;
        68: y = 16'b0111111101010011;
        69: y = 16'b0111111110010100;
        70: y = 16'b0111111111000101;
        71: y = 16'b0111111111101000;
        72: y = 16'b0111111111111011;
        73: y = 16'b0111111111111111;
        74: y = 16'b0111111111110011;
        75: y = 16'b0111111111011000;
        76: y = 16'b0111111110101110;
        77: y = 16'b0111111101110101;
        78: y = 16'b0111111100101101;
        79: y = 16'b0111111011010101;
        80: y = 16'b0111111001101110;
        81: y = 16'b0111110111111001;
        82: y = 16'b0111110101110100;
        83: y = 16'b0111110011100000;
        84: y = 16'b0111110000111101;
        85: y = 16'b0111101110001011;
        86: y = 16'b0111101011001011;
        87: y = 16'b0111100111111100;
        88: y = 16'b0111100100011111;
        89: y = 16'b0111100000110011;
        90: y = 16'b0111011100111000;
        91: y = 16'b0111011000110000;
        92: y = 16'b0111010100011001;
        93: y = 16'b0111001111110101;
        94: y = 16'b0111001011000010;
        95: y = 16'b0111000110000010;
        96: y = 16'b0111000000110100;
        97: y = 16'b0110111011011001;
        98: y = 16'b0110110101110001;
        99: y = 16'b0110101111111011;
        100: y = 16'b0110101001111001;
        101: y = 16'b0110100011101010;
        102: y = 16'b0110011101001111;
        103: y = 16'b0110010110100111;
        104: y = 16'b0110001111110011;
        105: y = 16'b0110001000110011;
        106: y = 16'b0110000001100111;
        107: y = 16'b0101111010010000;
        108: y = 16'b0101110010101110;
        109: y = 16'b0101101011000000;
        110: y = 16'b0101100011001000;
        111: y = 16'b0101011011000101;
        112: y = 16'b0101010010111000;
        113: y = 16'b0101001010100000;
        114: y = 16'b0101000001111111;
        115: y = 16'b0100111001010100;
        116: y = 16'b0100110000100000;
        117: y = 16'b0100100111100011;
        118: y = 16'b0100011110011101;
        119: y = 16'b0100010101001110;
        120: y = 16'b0100001011110111;
        121: y = 16'b0100000010011000;
        122: y = 16'b0011111000110010;
        123: y = 16'b0011101111000100;
        124: y = 16'b0011100101001111;
        125: y = 16'b0011011011010011;
        126: y = 16'b0011010001010000;
        127: y = 16'b0011000111000111;
        128: y = 16'b0010111100111001;
        129: y = 16'b0010110010100100;
        130: y = 16'b0010101000001011;
        131: y = 16'b0010011101101100;
        132: y = 16'b0010010011001001;
        133: y = 16'b0010001000100001;
        134: y = 16'b0001111101110101;
        135: y = 16'b0001110011000101;
        136: y = 16'b0001101000010010;
        137: y = 16'b0001011101011100;
        138: y = 16'b0001010010100011;
        139: y = 16'b0001000111101000;
        140: y = 16'b0000111100101010;
        141: y = 16'b0000110001101011;
        142: y = 16'b0000100110101010;
        143: y = 16'b0000011011101000;
        144: y = 16'b0000010000100101;
        145: y = 16'b0000000101100010;
        146: y = 16'b1111111010011110;
        147: y = 16'b1111101111011011;
        148: y = 16'b1111100100011000;
        149: y = 16'b1111011001010110;
        150: y = 16'b1111001110010101;
        151: y = 16'b1111000011010110;
        152: y = 16'b1110111000011000;
        153: y = 16'b1110101101011101;
        154: y = 16'b1110100010100100;
        155: y = 16'b1110010111101110;
        156: y = 16'b1110001100111011;
        157: y = 16'b1110000010001011;
        158: y = 16'b1101110111011111;
        159: y = 16'b1101101100110111;
        160: y = 16'b1101100010010100;
        161: y = 16'b1101010111110101;
        162: y = 16'b1101001101011100;
        163: y = 16'b1101000011000111;
        164: y = 16'b1100111000111001;
        165: y = 16'b1100101110110000;
        166: y = 16'b1100100100101101;
        167: y = 16'b1100011010110001;
        168: y = 16'b1100010000111100;
        169: y = 16'b1100000111001110;
        170: y = 16'b1011111101101000;
        171: y = 16'b1011110100001001;
        172: y = 16'b1011101010110010;
        173: y = 16'b1011100001100011;
        174: y = 16'b1011011000011101;
        175: y = 16'b1011001111100000;
        176: y = 16'b1011000110101100;
        177: y = 16'b1010111110000001;
        178: y = 16'b1010110101100000;
        179: y = 16'b1010101101001000;
        180: y = 16'b1010100100111011;
        181: y = 16'b1010011100111000;
        182: y = 16'b1010010101000000;
        183: y = 16'b1010001101010010;
        184: y = 16'b1010000101110000;
        185: y = 16'b1001111110011001;
        186: y = 16'b1001110111001101;
        187: y = 16'b1001110000001101;
        188: y = 16'b1001101001011001;
        189: y = 16'b1001100010110001;
        190: y = 16'b1001011100010110;
        191: y = 16'b1001010110000111;
        192: y = 16'b1001010000000101;
        193: y = 16'b1001001010001111;
        194: y = 16'b1001000100100111;
        195: y = 16'b1000111111001100;
        196: y = 16'b1000111001111110;
        197: y = 16'b1000110100111110;
        198: y = 16'b1000110000001011;
        199: y = 16'b1000101011100111;
        200: y = 16'b1000100111010000;
        201: y = 16'b1000100011001000;
        202: y = 16'b1000011111001101;
        203: y = 16'b1000011011100001;
        204: y = 16'b1000011000000100;
        205: y = 16'b1000010100110101;
        206: y = 16'b1000010001110101;
        207: y = 16'b1000001111000011;
        208: y = 16'b1000001100100000;
        209: y = 16'b1000001010001100;
        210: y = 16'b1000001000000111;
        211: y = 16'b1000000110010010;
        212: y = 16'b1000000100101011;
        213: y = 16'b1000000011010011;
        214: y = 16'b1000000010001011;
        215: y = 16'b1000000001010010;
        216: y = 16'b1000000000101000;
        217: y = 16'b1000000000001101;
        218: y = 16'b1000000000000001;
        219: y = 16'b1000000000000101;
        220: y = 16'b1000000000011000;
        221: y = 16'b1000000000111011;
        222: y = 16'b1000000001101100;
        223: y = 16'b1000000010101101;
        224: y = 16'b1000000011111101;
        225: y = 16'b1000000101011100;
        226: y = 16'b1000000111001011;
        227: y = 16'b1000001001001000;
        228: y = 16'b1000001011010100;
        229: y = 16'b1000001101110000;
        230: y = 16'b1000010000011010;
        231: y = 16'b1000010011010011;
        232: y = 16'b1000010110011010;
        233: y = 16'b1000011001110001;
        234: y = 16'b1000011101010110;
        235: y = 16'b1000100001001001;
        236: y = 16'b1000100101001010;
        237: y = 16'b1000101001011010;
        238: y = 16'b1000101101110111;
        239: y = 16'b1000110010100011;
        240: y = 16'b1000110111011100;
        241: y = 16'b1000111100100011;
        242: y = 16'b1001000001111000;
        243: y = 16'b1001000111011001;
        244: y = 16'b1001001101001000;
        245: y = 16'b1001010011000100;
        246: y = 16'b1001011001001101;
        247: y = 16'b1001011111100010;
        248: y = 16'b1001100110000100;
        249: y = 16'b1001101100110010;
        250: y = 16'b1001110011101100;
        251: y = 16'b1001111010110010;
        252: y = 16'b1010000010000011;
        253: y = 16'b1010001001100000;
        254: y = 16'b1010010001001000;
        255: y = 16'b1010011000111011;
        256: y = 16'b1010100000111000;
        257: y = 16'b1010101001000000;
        258: y = 16'b1010110001010011;
        259: y = 16'b1010111001101111;
        260: y = 16'b1011000010010101;
        261: y = 16'b1011001011000101;
        262: y = 16'b1011010011111101;
        263: y = 16'b1011011100111111;
        264: y = 16'b1011100110001001;
        265: y = 16'b1011101111011100;
        266: y = 16'b1011111000110111;
        267: y = 16'b1100000010011010;
        268: y = 16'b1100001100000100;
        269: y = 16'b1100010101110110;
        270: y = 16'b1100011111101110;
        271: y = 16'b1100101001101110;
        272: y = 16'b1100110011110011;
        273: y = 16'b1100111101111111;
        274: y = 16'b1101001000010001;
        275: y = 16'b1101010010101000;
        276: y = 16'b1101011101000100;
        277: y = 16'b1101100111100101;
        278: y = 16'b1101110010001011;
        279: y = 16'b1101111100110101;
        280: y = 16'b1110000111100011;
        281: y = 16'b1110010010010100;
        282: y = 16'b1110011101001001;
        283: y = 16'b1110101000000000;
        284: y = 16'b1110110010111010;
        285: y = 16'b1110111101110111;
        286: y = 16'b1111001000110101;
        287: y = 16'b1111010011110110;
        288: y = 16'b1111011110110111;
        289: y = 16'b1111101001111001;
        290: y = 16'b1111110100111101;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=349.23Hz, Fs=96000Hz, 16-bit

module lut_F
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 273;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001011101111;
        2: y = 16'b0000010111011110;
        3: y = 16'b0000100011001100;
        4: y = 16'b0000101110111001;
        5: y = 16'b0000111010100101;
        6: y = 16'b0001000110001110;
        7: y = 16'b0001010001110101;
        8: y = 16'b0001011101011001;
        9: y = 16'b0001101000111011;
        10: y = 16'b0001110100011000;
        11: y = 16'b0001111111110010;
        12: y = 16'b0010001011000111;
        13: y = 16'b0010010110011000;
        14: y = 16'b0010100001100100;
        15: y = 16'b0010101100101010;
        16: y = 16'b0010110111101010;
        17: y = 16'b0011000010100101;
        18: y = 16'b0011001101011000;
        19: y = 16'b0011011000000101;
        20: y = 16'b0011100010101011;
        21: y = 16'b0011101101001000;
        22: y = 16'b0011110111011110;
        23: y = 16'b0100000001101100;
        24: y = 16'b0100001011110001;
        25: y = 16'b0100010101101101;
        26: y = 16'b0100011111011111;
        27: y = 16'b0100101001001000;
        28: y = 16'b0100110010100111;
        29: y = 16'b0100111011111011;
        30: y = 16'b0101000101000101;
        31: y = 16'b0101001110000100;
        32: y = 16'b0101010110111000;
        33: y = 16'b0101011111100000;
        34: y = 16'b0101100111111101;
        35: y = 16'b0101110000001101;
        36: y = 16'b0101111000010001;
        37: y = 16'b0110000000001000;
        38: y = 16'b0110000111110010;
        39: y = 16'b0110001111001111;
        40: y = 16'b0110010110011111;
        41: y = 16'b0110011101100001;
        42: y = 16'b0110100100010101;
        43: y = 16'b0110101010111011;
        44: y = 16'b0110110001010010;
        45: y = 16'b0110110111011011;
        46: y = 16'b0110111101010101;
        47: y = 16'b0111000011000001;
        48: y = 16'b0111001000011101;
        49: y = 16'b0111001101101001;
        50: y = 16'b0111010010100110;
        51: y = 16'b0111010111010100;
        52: y = 16'b0111011011110001;
        53: y = 16'b0111011111111111;
        54: y = 16'b0111100011111100;
        55: y = 16'b0111100111101001;
        56: y = 16'b0111101011000110;
        57: y = 16'b0111101110010010;
        58: y = 16'b0111110001001110;
        59: y = 16'b0111110011111001;
        60: y = 16'b0111110110010011;
        61: y = 16'b0111111000011100;
        62: y = 16'b0111111010010100;
        63: y = 16'b0111111011111011;
        64: y = 16'b0111111101010001;
        65: y = 16'b0111111110010110;
        66: y = 16'b0111111111001001;
        67: y = 16'b0111111111101100;
        68: y = 16'b0111111111111101;
        69: y = 16'b0111111111111101;
        70: y = 16'b0111111111101100;
        71: y = 16'b0111111111001001;
        72: y = 16'b0111111110010110;
        73: y = 16'b0111111101010001;
        74: y = 16'b0111111011111011;
        75: y = 16'b0111111010010100;
        76: y = 16'b0111111000011100;
        77: y = 16'b0111110110010011;
        78: y = 16'b0111110011111001;
        79: y = 16'b0111110001001110;
        80: y = 16'b0111101110010010;
        81: y = 16'b0111101011000110;
        82: y = 16'b0111100111101001;
        83: y = 16'b0111100011111100;
        84: y = 16'b0111011111111111;
        85: y = 16'b0111011011110001;
        86: y = 16'b0111010111010100;
        87: y = 16'b0111010010100110;
        88: y = 16'b0111001101101001;
        89: y = 16'b0111001000011101;
        90: y = 16'b0111000011000001;
        91: y = 16'b0110111101010101;
        92: y = 16'b0110110111011011;
        93: y = 16'b0110110001010010;
        94: y = 16'b0110101010111011;
        95: y = 16'b0110100100010101;
        96: y = 16'b0110011101100001;
        97: y = 16'b0110010110011111;
        98: y = 16'b0110001111001111;
        99: y = 16'b0110000111110010;
        100: y = 16'b0110000000001000;
        101: y = 16'b0101111000010001;
        102: y = 16'b0101110000001101;
        103: y = 16'b0101100111111101;
        104: y = 16'b0101011111100000;
        105: y = 16'b0101010110111000;
        106: y = 16'b0101001110000100;
        107: y = 16'b0101000101000101;
        108: y = 16'b0100111011111011;
        109: y = 16'b0100110010100111;
        110: y = 16'b0100101001001000;
        111: y = 16'b0100011111011111;
        112: y = 16'b0100010101101101;
        113: y = 16'b0100001011110001;
        114: y = 16'b0100000001101100;
        115: y = 16'b0011110111011110;
        116: y = 16'b0011101101001000;
        117: y = 16'b0011100010101011;
        118: y = 16'b0011011000000101;
        119: y = 16'b0011001101011000;
        120: y = 16'b0011000010100101;
        121: y = 16'b0010110111101010;
        122: y = 16'b0010101100101010;
        123: y = 16'b0010100001100100;
        124: y = 16'b0010010110011000;
        125: y = 16'b0010001011000111;
        126: y = 16'b0001111111110010;
        127: y = 16'b0001110100011000;
        128: y = 16'b0001101000111011;
        129: y = 16'b0001011101011001;
        130: y = 16'b0001010001110101;
        131: y = 16'b0001000110001110;
        132: y = 16'b0000111010100101;
        133: y = 16'b0000101110111001;
        134: y = 16'b0000100011001100;
        135: y = 16'b0000010111011110;
        136: y = 16'b0000001011101111;
        137: y = 16'b0000000000000000;
        138: y = 16'b1111110100010001;
        139: y = 16'b1111101000100010;
        140: y = 16'b1111011100110100;
        141: y = 16'b1111010001000111;
        142: y = 16'b1111000101011011;
        143: y = 16'b1110111001110010;
        144: y = 16'b1110101110001011;
        145: y = 16'b1110100010100111;
        146: y = 16'b1110010111000101;
        147: y = 16'b1110001011101000;
        148: y = 16'b1110000000001110;
        149: y = 16'b1101110100111001;
        150: y = 16'b1101101001101000;
        151: y = 16'b1101011110011100;
        152: y = 16'b1101010011010110;
        153: y = 16'b1101001000010110;
        154: y = 16'b1100111101011011;
        155: y = 16'b1100110010101000;
        156: y = 16'b1100100111111011;
        157: y = 16'b1100011101010101;
        158: y = 16'b1100010010111000;
        159: y = 16'b1100001000100010;
        160: y = 16'b1011111110010100;
        161: y = 16'b1011110100001111;
        162: y = 16'b1011101010010011;
        163: y = 16'b1011100000100001;
        164: y = 16'b1011010110111000;
        165: y = 16'b1011001101011001;
        166: y = 16'b1011000100000101;
        167: y = 16'b1010111010111011;
        168: y = 16'b1010110001111100;
        169: y = 16'b1010101001001000;
        170: y = 16'b1010100000100000;
        171: y = 16'b1010011000000011;
        172: y = 16'b1010001111110011;
        173: y = 16'b1010000111101111;
        174: y = 16'b1001111111111000;
        175: y = 16'b1001111000001110;
        176: y = 16'b1001110000110001;
        177: y = 16'b1001101001100001;
        178: y = 16'b1001100010011111;
        179: y = 16'b1001011011101011;
        180: y = 16'b1001010101000101;
        181: y = 16'b1001001110101110;
        182: y = 16'b1001001000100101;
        183: y = 16'b1001000010101011;
        184: y = 16'b1000111100111111;
        185: y = 16'b1000110111100011;
        186: y = 16'b1000110010010111;
        187: y = 16'b1000101101011010;
        188: y = 16'b1000101000101100;
        189: y = 16'b1000100100001111;
        190: y = 16'b1000100000000001;
        191: y = 16'b1000011100000100;
        192: y = 16'b1000011000010111;
        193: y = 16'b1000010100111010;
        194: y = 16'b1000010001101110;
        195: y = 16'b1000001110110010;
        196: y = 16'b1000001100000111;
        197: y = 16'b1000001001101101;
        198: y = 16'b1000000111100100;
        199: y = 16'b1000000101101100;
        200: y = 16'b1000000100000101;
        201: y = 16'b1000000010101111;
        202: y = 16'b1000000001101010;
        203: y = 16'b1000000000110111;
        204: y = 16'b1000000000010100;
        205: y = 16'b1000000000000011;
        206: y = 16'b1000000000000011;
        207: y = 16'b1000000000010100;
        208: y = 16'b1000000000110111;
        209: y = 16'b1000000001101010;
        210: y = 16'b1000000010101111;
        211: y = 16'b1000000100000101;
        212: y = 16'b1000000101101100;
        213: y = 16'b1000000111100100;
        214: y = 16'b1000001001101101;
        215: y = 16'b1000001100000111;
        216: y = 16'b1000001110110010;
        217: y = 16'b1000010001101110;
        218: y = 16'b1000010100111010;
        219: y = 16'b1000011000010111;
        220: y = 16'b1000011100000100;
        221: y = 16'b1000100000000001;
        222: y = 16'b1000100100001111;
        223: y = 16'b1000101000101100;
        224: y = 16'b1000101101011010;
        225: y = 16'b1000110010010111;
        226: y = 16'b1000110111100011;
        227: y = 16'b1000111100111111;
        228: y = 16'b1001000010101011;
        229: y = 16'b1001001000100101;
        230: y = 16'b1001001110101110;
        231: y = 16'b1001010101000101;
        232: y = 16'b1001011011101011;
        233: y = 16'b1001100010011111;
        234: y = 16'b1001101001100001;
        235: y = 16'b1001110000110001;
        236: y = 16'b1001111000001110;
        237: y = 16'b1001111111111000;
        238: y = 16'b1010000111101111;
        239: y = 16'b1010001111110011;
        240: y = 16'b1010011000000011;
        241: y = 16'b1010100000100000;
        242: y = 16'b1010101001001000;
        243: y = 16'b1010110001111100;
        244: y = 16'b1010111010111011;
        245: y = 16'b1011000100000101;
        246: y = 16'b1011001101011001;
        247: y = 16'b1011010110111000;
        248: y = 16'b1011100000100001;
        249: y = 16'b1011101010010011;
        250: y = 16'b1011110100001111;
        251: y = 16'b1011111110010100;
        252: y = 16'b1100001000100010;
        253: y = 16'b1100010010111000;
        254: y = 16'b1100011101010101;
        255: y = 16'b1100100111111011;
        256: y = 16'b1100110010101000;
        257: y = 16'b1100111101011011;
        258: y = 16'b1101001000010110;
        259: y = 16'b1101010011010110;
        260: y = 16'b1101011110011100;
        261: y = 16'b1101101001101000;
        262: y = 16'b1101110100111001;
        263: y = 16'b1110000000001110;
        264: y = 16'b1110001011101000;
        265: y = 16'b1110010111000101;
        266: y = 16'b1110100010100111;
        267: y = 16'b1110101110001011;
        268: y = 16'b1110111001110010;
        269: y = 16'b1111000101011011;
        270: y = 16'b1111010001000111;
        271: y = 16'b1111011100110100;
        272: y = 16'b1111101000100010;
        273: y = 16'b1111110100010001;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=369.99Hz, Fs=96000Hz, 16-bit

module lut_Fs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 258;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001100011011;
        2: y = 16'b0000011000110101;
        3: y = 16'b0000100101001111;
        4: y = 16'b0000110001100111;
        5: y = 16'b0000111101111101;
        6: y = 16'b0001001010010001;
        7: y = 16'b0001010110100010;
        8: y = 16'b0001100010101111;
        9: y = 16'b0001101110111001;
        10: y = 16'b0001111010111111;
        11: y = 16'b0010000111000001;
        12: y = 16'b0010010010111101;
        13: y = 16'b0010011110110011;
        14: y = 16'b0010101010100100;
        15: y = 16'b0010110110001110;
        16: y = 16'b0011000001110010;
        17: y = 16'b0011001101001110;
        18: y = 16'b0011011000100010;
        19: y = 16'b0011100011101110;
        20: y = 16'b0011101110110010;
        21: y = 16'b0011111001101100;
        22: y = 16'b0100000100011101;
        23: y = 16'b0100001111000101;
        24: y = 16'b0100011001100010;
        25: y = 16'b0100100011110101;
        26: y = 16'b0100101101111100;
        27: y = 16'b0100110111111000;
        28: y = 16'b0101000001101001;
        29: y = 16'b0101001011001101;
        30: y = 16'b0101010100100101;
        31: y = 16'b0101011101110000;
        32: y = 16'b0101100110101110;
        33: y = 16'b0101101111011110;
        34: y = 16'b0101111000000001;
        35: y = 16'b0110000000010101;
        36: y = 16'b0110001000011011;
        37: y = 16'b0110010000010010;
        38: y = 16'b0110010111111010;
        39: y = 16'b0110011111010011;
        40: y = 16'b0110100110011100;
        41: y = 16'b0110101101010101;
        42: y = 16'b0110110011111110;
        43: y = 16'b0110111010010111;
        44: y = 16'b0111000000011110;
        45: y = 16'b0111000110010101;
        46: y = 16'b0111001011111011;
        47: y = 16'b0111010001010000;
        48: y = 16'b0111010110010011;
        49: y = 16'b0111011011000100;
        50: y = 16'b0111011111100100;
        51: y = 16'b0111100011110001;
        52: y = 16'b0111100111101100;
        53: y = 16'b0111101011010101;
        54: y = 16'b0111101110101011;
        55: y = 16'b0111110001101111;
        56: y = 16'b0111110100100000;
        57: y = 16'b0111110110111110;
        58: y = 16'b0111111001001001;
        59: y = 16'b0111111011000001;
        60: y = 16'b0111111100100110;
        61: y = 16'b0111111101111000;
        62: y = 16'b0111111110110110;
        63: y = 16'b0111111111100001;
        64: y = 16'b0111111111111010;
        65: y = 16'b0111111111111110;
        66: y = 16'b0111111111110000;
        67: y = 16'b0111111111001110;
        68: y = 16'b0111111110011001;
        69: y = 16'b0111111101010001;
        70: y = 16'b0111111011110110;
        71: y = 16'b0111111010000111;
        72: y = 16'b0111111000000101;
        73: y = 16'b0111110101110001;
        74: y = 16'b0111110011001001;
        75: y = 16'b0111110000001111;
        76: y = 16'b0111101101000010;
        77: y = 16'b0111101001100011;
        78: y = 16'b0111100101110001;
        79: y = 16'b0111100001101100;
        80: y = 16'b0111011101010110;
        81: y = 16'b0111011000101110;
        82: y = 16'b0111010011110100;
        83: y = 16'b0111001110101000;
        84: y = 16'b0111001001001011;
        85: y = 16'b0111000011011100;
        86: y = 16'b0110111101011101;
        87: y = 16'b0110110111001100;
        88: y = 16'b0110110000101100;
        89: y = 16'b0110101001111011;
        90: y = 16'b0110100010111001;
        91: y = 16'b0110011011101001;
        92: y = 16'b0110010100001000;
        93: y = 16'b0110001100011001;
        94: y = 16'b0110000100011010;
        95: y = 16'b0101111100001101;
        96: y = 16'b0101110011110001;
        97: y = 16'b0101101011001000;
        98: y = 16'b0101100010010001;
        99: y = 16'b0101011001001100;
        100: y = 16'b0101001111111011;
        101: y = 16'b0101000110011101;
        102: y = 16'b0100111100110010;
        103: y = 16'b0100110010111100;
        104: y = 16'b0100101000111010;
        105: y = 16'b0100011110101101;
        106: y = 16'b0100010100010101;
        107: y = 16'b0100001001110010;
        108: y = 16'b0011111111000110;
        109: y = 16'b0011110100010000;
        110: y = 16'b0011101001010001;
        111: y = 16'b0011011110001001;
        112: y = 16'b0011010010111001;
        113: y = 16'b0011000111100001;
        114: y = 16'b0010111100000001;
        115: y = 16'b0010110000011010;
        116: y = 16'b0010100100101100;
        117: y = 16'b0010011000111001;
        118: y = 16'b0010001100111111;
        119: y = 16'b0010000001000001;
        120: y = 16'b0001110100111101;
        121: y = 16'b0001101000110101;
        122: y = 16'b0001011100101001;
        123: y = 16'b0001010000011010;
        124: y = 16'b0001000100000111;
        125: y = 16'b0000110111110010;
        126: y = 16'b0000101011011011;
        127: y = 16'b0000011111000010;
        128: y = 16'b0000010010101000;
        129: y = 16'b0000000110001101;
        130: y = 16'b1111111001110011;
        131: y = 16'b1111101101011000;
        132: y = 16'b1111100000111110;
        133: y = 16'b1111010100100101;
        134: y = 16'b1111001000001110;
        135: y = 16'b1110111011111001;
        136: y = 16'b1110101111100110;
        137: y = 16'b1110100011010111;
        138: y = 16'b1110010111001011;
        139: y = 16'b1110001011000011;
        140: y = 16'b1101111110111111;
        141: y = 16'b1101110011000001;
        142: y = 16'b1101100111000111;
        143: y = 16'b1101011011010100;
        144: y = 16'b1101001111100110;
        145: y = 16'b1101000011111111;
        146: y = 16'b1100111000011111;
        147: y = 16'b1100101101000111;
        148: y = 16'b1100100001110111;
        149: y = 16'b1100010110101111;
        150: y = 16'b1100001011110000;
        151: y = 16'b1100000000111010;
        152: y = 16'b1011110110001110;
        153: y = 16'b1011101011101011;
        154: y = 16'b1011100001010011;
        155: y = 16'b1011010111000110;
        156: y = 16'b1011001101000100;
        157: y = 16'b1011000011001110;
        158: y = 16'b1010111001100011;
        159: y = 16'b1010110000000101;
        160: y = 16'b1010100110110100;
        161: y = 16'b1010011101101111;
        162: y = 16'b1010010100111000;
        163: y = 16'b1010001100001111;
        164: y = 16'b1010000011110011;
        165: y = 16'b1001111011100110;
        166: y = 16'b1001110011100111;
        167: y = 16'b1001101011111000;
        168: y = 16'b1001100100010111;
        169: y = 16'b1001011101000111;
        170: y = 16'b1001010110000101;
        171: y = 16'b1001001111010100;
        172: y = 16'b1001001000110100;
        173: y = 16'b1001000010100011;
        174: y = 16'b1000111100100100;
        175: y = 16'b1000110110110101;
        176: y = 16'b1000110001011000;
        177: y = 16'b1000101100001100;
        178: y = 16'b1000100111010010;
        179: y = 16'b1000100010101010;
        180: y = 16'b1000011110010100;
        181: y = 16'b1000011010001111;
        182: y = 16'b1000010110011101;
        183: y = 16'b1000010010111110;
        184: y = 16'b1000001111110001;
        185: y = 16'b1000001100110111;
        186: y = 16'b1000001010001111;
        187: y = 16'b1000000111111011;
        188: y = 16'b1000000101111001;
        189: y = 16'b1000000100001010;
        190: y = 16'b1000000010101111;
        191: y = 16'b1000000001100111;
        192: y = 16'b1000000000110010;
        193: y = 16'b1000000000010000;
        194: y = 16'b1000000000000010;
        195: y = 16'b1000000000000110;
        196: y = 16'b1000000000011111;
        197: y = 16'b1000000001001010;
        198: y = 16'b1000000010001000;
        199: y = 16'b1000000011011010;
        200: y = 16'b1000000100111111;
        201: y = 16'b1000000110110111;
        202: y = 16'b1000001001000010;
        203: y = 16'b1000001011100000;
        204: y = 16'b1000001110010001;
        205: y = 16'b1000010001010101;
        206: y = 16'b1000010100101011;
        207: y = 16'b1000011000010100;
        208: y = 16'b1000011100001111;
        209: y = 16'b1000100000011100;
        210: y = 16'b1000100100111100;
        211: y = 16'b1000101001101101;
        212: y = 16'b1000101110110000;
        213: y = 16'b1000110100000101;
        214: y = 16'b1000111001101011;
        215: y = 16'b1000111111100010;
        216: y = 16'b1001000101101001;
        217: y = 16'b1001001100000010;
        218: y = 16'b1001010010101011;
        219: y = 16'b1001011001100100;
        220: y = 16'b1001100000101101;
        221: y = 16'b1001101000000110;
        222: y = 16'b1001101111101110;
        223: y = 16'b1001110111100101;
        224: y = 16'b1001111111101011;
        225: y = 16'b1010000111111111;
        226: y = 16'b1010010000100010;
        227: y = 16'b1010011001010010;
        228: y = 16'b1010100010010000;
        229: y = 16'b1010101011011011;
        230: y = 16'b1010110100110011;
        231: y = 16'b1010111110010111;
        232: y = 16'b1011001000001000;
        233: y = 16'b1011010010000100;
        234: y = 16'b1011011100001011;
        235: y = 16'b1011100110011110;
        236: y = 16'b1011110000111011;
        237: y = 16'b1011111011100011;
        238: y = 16'b1100000110010100;
        239: y = 16'b1100010001001110;
        240: y = 16'b1100011100010010;
        241: y = 16'b1100100111011110;
        242: y = 16'b1100110010110010;
        243: y = 16'b1100111110001110;
        244: y = 16'b1101001001110010;
        245: y = 16'b1101010101011100;
        246: y = 16'b1101100001001101;
        247: y = 16'b1101101101000011;
        248: y = 16'b1101111000111111;
        249: y = 16'b1110000101000001;
        250: y = 16'b1110010001000111;
        251: y = 16'b1110011101010001;
        252: y = 16'b1110101001011110;
        253: y = 16'b1110110101101111;
        254: y = 16'b1111000010000011;
        255: y = 16'b1111001110011001;
        256: y = 16'b1111011010110001;
        257: y = 16'b1111100111001011;
        258: y = 16'b1111110011100101;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=392.0Hz, Fs=96000Hz, 16-bit

module lut_G
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 243;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001101001100;
        2: y = 16'b0000011010010111;
        3: y = 16'b0000100111100001;
        4: y = 16'b0000110100101001;
        5: y = 16'b0001000001101111;
        6: y = 16'b0001001110110011;
        7: y = 16'b0001011011110010;
        8: y = 16'b0001101000101111;
        9: y = 16'b0001110101100110;
        10: y = 16'b0010000010011001;
        11: y = 16'b0010001111000110;
        12: y = 16'b0010011011101101;
        13: y = 16'b0010101000001101;
        14: y = 16'b0010110100100111;
        15: y = 16'b0011000000111000;
        16: y = 16'b0011001101000010;
        17: y = 16'b0011011001000010;
        18: y = 16'b0011100100111010;
        19: y = 16'b0011110000101000;
        20: y = 16'b0011111100001011;
        21: y = 16'b0100000111100100;
        22: y = 16'b0100010010110010;
        23: y = 16'b0100011101110100;
        24: y = 16'b0100101000101010;
        25: y = 16'b0100110011010011;
        26: y = 16'b0100111101110000;
        27: y = 16'b0101000111111110;
        28: y = 16'b0101010001111111;
        29: y = 16'b0101011011110010;
        30: y = 16'b0101100101010110;
        31: y = 16'b0101101110101010;
        32: y = 16'b0101110111101111;
        33: y = 16'b0110000000100100;
        34: y = 16'b0110001001001001;
        35: y = 16'b0110010001011101;
        36: y = 16'b0110011001100000;
        37: y = 16'b0110100001010010;
        38: y = 16'b0110101000110010;
        39: y = 16'b0110110000000000;
        40: y = 16'b0110110110111100;
        41: y = 16'b0110111101100101;
        42: y = 16'b0111000011111011;
        43: y = 16'b0111001001111110;
        44: y = 16'b0111001111101101;
        45: y = 16'b0111010101001001;
        46: y = 16'b0111011010010001;
        47: y = 16'b0111011111000101;
        48: y = 16'b0111100011100100;
        49: y = 16'b0111100111101111;
        50: y = 16'b0111101011100101;
        51: y = 16'b0111101111000111;
        52: y = 16'b0111110010010011;
        53: y = 16'b0111110101001010;
        54: y = 16'b0111110111101100;
        55: y = 16'b0111111001111001;
        56: y = 16'b0111111011110000;
        57: y = 16'b0111111101010001;
        58: y = 16'b0111111110011101;
        59: y = 16'b0111111111010100;
        60: y = 16'b0111111111110100;
        61: y = 16'b0111111111111111;
        62: y = 16'b0111111111110100;
        63: y = 16'b0111111111010100;
        64: y = 16'b0111111110011101;
        65: y = 16'b0111111101010001;
        66: y = 16'b0111111011110000;
        67: y = 16'b0111111001111001;
        68: y = 16'b0111110111101100;
        69: y = 16'b0111110101001010;
        70: y = 16'b0111110010010011;
        71: y = 16'b0111101111000111;
        72: y = 16'b0111101011100101;
        73: y = 16'b0111100111101111;
        74: y = 16'b0111100011100100;
        75: y = 16'b0111011111000101;
        76: y = 16'b0111011010010001;
        77: y = 16'b0111010101001001;
        78: y = 16'b0111001111101101;
        79: y = 16'b0111001001111110;
        80: y = 16'b0111000011111011;
        81: y = 16'b0110111101100101;
        82: y = 16'b0110110110111100;
        83: y = 16'b0110110000000000;
        84: y = 16'b0110101000110010;
        85: y = 16'b0110100001010010;
        86: y = 16'b0110011001100000;
        87: y = 16'b0110010001011101;
        88: y = 16'b0110001001001001;
        89: y = 16'b0110000000100100;
        90: y = 16'b0101110111101111;
        91: y = 16'b0101101110101010;
        92: y = 16'b0101100101010110;
        93: y = 16'b0101011011110010;
        94: y = 16'b0101010001111111;
        95: y = 16'b0101000111111110;
        96: y = 16'b0100111101110000;
        97: y = 16'b0100110011010011;
        98: y = 16'b0100101000101010;
        99: y = 16'b0100011101110100;
        100: y = 16'b0100010010110010;
        101: y = 16'b0100000111100100;
        102: y = 16'b0011111100001011;
        103: y = 16'b0011110000101000;
        104: y = 16'b0011100100111010;
        105: y = 16'b0011011001000010;
        106: y = 16'b0011001101000010;
        107: y = 16'b0011000000111000;
        108: y = 16'b0010110100100111;
        109: y = 16'b0010101000001101;
        110: y = 16'b0010011011101101;
        111: y = 16'b0010001111000110;
        112: y = 16'b0010000010011001;
        113: y = 16'b0001110101100110;
        114: y = 16'b0001101000101111;
        115: y = 16'b0001011011110010;
        116: y = 16'b0001001110110011;
        117: y = 16'b0001000001101111;
        118: y = 16'b0000110100101001;
        119: y = 16'b0000100111100001;
        120: y = 16'b0000011010010111;
        121: y = 16'b0000001101001100;
        122: y = 16'b0000000000000000;
        123: y = 16'b1111110010110100;
        124: y = 16'b1111100101101001;
        125: y = 16'b1111011000011111;
        126: y = 16'b1111001011010111;
        127: y = 16'b1110111110010001;
        128: y = 16'b1110110001001101;
        129: y = 16'b1110100100001110;
        130: y = 16'b1110010111010001;
        131: y = 16'b1110001010011010;
        132: y = 16'b1101111101100111;
        133: y = 16'b1101110000111010;
        134: y = 16'b1101100100010011;
        135: y = 16'b1101010111110011;
        136: y = 16'b1101001011011001;
        137: y = 16'b1100111111001000;
        138: y = 16'b1100110010111110;
        139: y = 16'b1100100110111110;
        140: y = 16'b1100011011000110;
        141: y = 16'b1100001111011000;
        142: y = 16'b1100000011110101;
        143: y = 16'b1011111000011100;
        144: y = 16'b1011101101001110;
        145: y = 16'b1011100010001100;
        146: y = 16'b1011010111010110;
        147: y = 16'b1011001100101101;
        148: y = 16'b1011000010010000;
        149: y = 16'b1010111000000010;
        150: y = 16'b1010101110000001;
        151: y = 16'b1010100100001110;
        152: y = 16'b1010011010101010;
        153: y = 16'b1010010001010110;
        154: y = 16'b1010001000010001;
        155: y = 16'b1001111111011100;
        156: y = 16'b1001110110110111;
        157: y = 16'b1001101110100011;
        158: y = 16'b1001100110100000;
        159: y = 16'b1001011110101110;
        160: y = 16'b1001010111001110;
        161: y = 16'b1001010000000000;
        162: y = 16'b1001001001000100;
        163: y = 16'b1001000010011011;
        164: y = 16'b1000111100000101;
        165: y = 16'b1000110110000010;
        166: y = 16'b1000110000010011;
        167: y = 16'b1000101010110111;
        168: y = 16'b1000100101101111;
        169: y = 16'b1000100000111011;
        170: y = 16'b1000011100011100;
        171: y = 16'b1000011000010001;
        172: y = 16'b1000010100011011;
        173: y = 16'b1000010000111001;
        174: y = 16'b1000001101101101;
        175: y = 16'b1000001010110110;
        176: y = 16'b1000001000010100;
        177: y = 16'b1000000110000111;
        178: y = 16'b1000000100010000;
        179: y = 16'b1000000010101111;
        180: y = 16'b1000000001100011;
        181: y = 16'b1000000000101100;
        182: y = 16'b1000000000001100;
        183: y = 16'b1000000000000001;
        184: y = 16'b1000000000001100;
        185: y = 16'b1000000000101100;
        186: y = 16'b1000000001100011;
        187: y = 16'b1000000010101111;
        188: y = 16'b1000000100010000;
        189: y = 16'b1000000110000111;
        190: y = 16'b1000001000010100;
        191: y = 16'b1000001010110110;
        192: y = 16'b1000001101101101;
        193: y = 16'b1000010000111001;
        194: y = 16'b1000010100011011;
        195: y = 16'b1000011000010001;
        196: y = 16'b1000011100011100;
        197: y = 16'b1000100000111011;
        198: y = 16'b1000100101101111;
        199: y = 16'b1000101010110111;
        200: y = 16'b1000110000010011;
        201: y = 16'b1000110110000010;
        202: y = 16'b1000111100000101;
        203: y = 16'b1001000010011011;
        204: y = 16'b1001001001000100;
        205: y = 16'b1001010000000000;
        206: y = 16'b1001010111001110;
        207: y = 16'b1001011110101110;
        208: y = 16'b1001100110100000;
        209: y = 16'b1001101110100011;
        210: y = 16'b1001110110110111;
        211: y = 16'b1001111111011100;
        212: y = 16'b1010001000010001;
        213: y = 16'b1010010001010110;
        214: y = 16'b1010011010101010;
        215: y = 16'b1010100100001110;
        216: y = 16'b1010101110000001;
        217: y = 16'b1010111000000010;
        218: y = 16'b1011000010010000;
        219: y = 16'b1011001100101101;
        220: y = 16'b1011010111010110;
        221: y = 16'b1011100010001100;
        222: y = 16'b1011101101001110;
        223: y = 16'b1011111000011100;
        224: y = 16'b1100000011110101;
        225: y = 16'b1100001111011000;
        226: y = 16'b1100011011000110;
        227: y = 16'b1100100110111110;
        228: y = 16'b1100110010111110;
        229: y = 16'b1100111111001000;
        230: y = 16'b1101001011011001;
        231: y = 16'b1101010111110011;
        232: y = 16'b1101100100010011;
        233: y = 16'b1101110000111010;
        234: y = 16'b1101111101100111;
        235: y = 16'b1110001010011010;
        236: y = 16'b1110010111010001;
        237: y = 16'b1110100100001110;
        238: y = 16'b1110110001001101;
        239: y = 16'b1110111110010001;
        240: y = 16'b1111001011010111;
        241: y = 16'b1111011000011111;
        242: y = 16'b1111100101101001;
        243: y = 16'b1111110010110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=415.3Hz, Fs=96000Hz, 16-bit

module lut_Gs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 230;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001101111011;
        2: y = 16'b0000011011110110;
        3: y = 16'b0000101001101111;
        4: y = 16'b0000110111100110;
        5: y = 16'b0001000101011011;
        6: y = 16'b0001010011001100;
        7: y = 16'b0001100000111001;
        8: y = 16'b0001101110100010;
        9: y = 16'b0001111100000101;
        10: y = 16'b0010001001100011;
        11: y = 16'b0010010110111010;
        12: y = 16'b0010100100001010;
        13: y = 16'b0010110001010010;
        14: y = 16'b0010111110010010;
        15: y = 16'b0011001011001001;
        16: y = 16'b0011010111110110;
        17: y = 16'b0011100100011001;
        18: y = 16'b0011110000110001;
        19: y = 16'b0011111100111110;
        20: y = 16'b0100001000111111;
        21: y = 16'b0100010100110011;
        22: y = 16'b0100100000011010;
        23: y = 16'b0100101011110100;
        24: y = 16'b0100110110111111;
        25: y = 16'b0101000001111100;
        26: y = 16'b0101001100101001;
        27: y = 16'b0101010111000110;
        28: y = 16'b0101100001010100;
        29: y = 16'b0101101011010000;
        30: y = 16'b0101110100111100;
        31: y = 16'b0101111110010110;
        32: y = 16'b0110000111011101;
        33: y = 16'b0110010000010010;
        34: y = 16'b0110011000110100;
        35: y = 16'b0110100001000011;
        36: y = 16'b0110101000111110;
        37: y = 16'b0110110000100101;
        38: y = 16'b0110110111111000;
        39: y = 16'b0110111110110101;
        40: y = 16'b0111000101011110;
        41: y = 16'b0111001011110001;
        42: y = 16'b0111010001101110;
        43: y = 16'b0111010111010101;
        44: y = 16'b0111011100100110;
        45: y = 16'b0111100001100000;
        46: y = 16'b0111100110000100;
        47: y = 16'b0111101010010000;
        48: y = 16'b0111101110000101;
        49: y = 16'b0111110001100011;
        50: y = 16'b0111110100101010;
        51: y = 16'b0111110111011000;
        52: y = 16'b0111111001101111;
        53: y = 16'b0111111011101110;
        54: y = 16'b0111111101010101;
        55: y = 16'b0111111110100011;
        56: y = 16'b0111111111011010;
        57: y = 16'b0111111111111000;
        58: y = 16'b0111111111111110;
        59: y = 16'b0111111111101100;
        60: y = 16'b0111111111000010;
        61: y = 16'b0111111101111111;
        62: y = 16'b0111111100100100;
        63: y = 16'b0111111010110001;
        64: y = 16'b0111111000100111;
        65: y = 16'b0111110110000100;
        66: y = 16'b0111110011001001;
        67: y = 16'b0111101111110111;
        68: y = 16'b0111101100001110;
        69: y = 16'b0111101000001101;
        70: y = 16'b0111100011110101;
        71: y = 16'b0111011111000110;
        72: y = 16'b0111011010000000;
        73: y = 16'b0111010100100100;
        74: y = 16'b0111001110110010;
        75: y = 16'b0111001000101010;
        76: y = 16'b0111000010001100;
        77: y = 16'b0110111011011001;
        78: y = 16'b0110110100010001;
        79: y = 16'b0110101100110100;
        80: y = 16'b0110100101000011;
        81: y = 16'b0110011100111110;
        82: y = 16'b0110010100100110;
        83: y = 16'b0110001011111010;
        84: y = 16'b0110000010111100;
        85: y = 16'b0101111001101011;
        86: y = 16'b0101110000001000;
        87: y = 16'b0101100110010100;
        88: y = 16'b0101011100001111;
        89: y = 16'b0101010001111010;
        90: y = 16'b0101000111010100;
        91: y = 16'b0100111100011111;
        92: y = 16'b0100110001011011;
        93: y = 16'b0100100110001001;
        94: y = 16'b0100011010101000;
        95: y = 16'b0100001110111011;
        96: y = 16'b0100000011000000;
        97: y = 16'b0011110110111001;
        98: y = 16'b0011101010100111;
        99: y = 16'b0011011110001001;
        100: y = 16'b0011010001100001;
        101: y = 16'b0011000100101111;
        102: y = 16'b0010110111110011;
        103: y = 16'b0010101010101111;
        104: y = 16'b0010011101100011;
        105: y = 16'b0010010000010000;
        106: y = 16'b0010000010110101;
        107: y = 16'b0001110101010100;
        108: y = 16'b0001100111101110;
        109: y = 16'b0001011010000011;
        110: y = 16'b0001001100010100;
        111: y = 16'b0000111110100001;
        112: y = 16'b0000110000101011;
        113: y = 16'b0000100010110010;
        114: y = 16'b0000010100111001;
        115: y = 16'b0000000110111110;
        116: y = 16'b1111111001000010;
        117: y = 16'b1111101011000111;
        118: y = 16'b1111011101001110;
        119: y = 16'b1111001111010101;
        120: y = 16'b1111000001011111;
        121: y = 16'b1110110011101100;
        122: y = 16'b1110100101111101;
        123: y = 16'b1110011000010010;
        124: y = 16'b1110001010101100;
        125: y = 16'b1101111101001011;
        126: y = 16'b1101101111110000;
        127: y = 16'b1101100010011101;
        128: y = 16'b1101010101010001;
        129: y = 16'b1101001000001101;
        130: y = 16'b1100111011010001;
        131: y = 16'b1100101110011111;
        132: y = 16'b1100100001110111;
        133: y = 16'b1100010101011001;
        134: y = 16'b1100001001000111;
        135: y = 16'b1011111101000000;
        136: y = 16'b1011110001000101;
        137: y = 16'b1011100101011000;
        138: y = 16'b1011011001110111;
        139: y = 16'b1011001110100101;
        140: y = 16'b1011000011100001;
        141: y = 16'b1010111000101100;
        142: y = 16'b1010101110000110;
        143: y = 16'b1010100011110001;
        144: y = 16'b1010011001101100;
        145: y = 16'b1010001111111000;
        146: y = 16'b1010000110010101;
        147: y = 16'b1001111101000100;
        148: y = 16'b1001110100000110;
        149: y = 16'b1001101011011010;
        150: y = 16'b1001100011000010;
        151: y = 16'b1001011010111101;
        152: y = 16'b1001010011001100;
        153: y = 16'b1001001011101111;
        154: y = 16'b1001000100100111;
        155: y = 16'b1000111101110100;
        156: y = 16'b1000110111010110;
        157: y = 16'b1000110001001110;
        158: y = 16'b1000101011011100;
        159: y = 16'b1000100110000000;
        160: y = 16'b1000100000111010;
        161: y = 16'b1000011100001011;
        162: y = 16'b1000010111110011;
        163: y = 16'b1000010011110010;
        164: y = 16'b1000010000001001;
        165: y = 16'b1000001100110111;
        166: y = 16'b1000001001111100;
        167: y = 16'b1000000111011001;
        168: y = 16'b1000000101001111;
        169: y = 16'b1000000011011100;
        170: y = 16'b1000000010000001;
        171: y = 16'b1000000000111110;
        172: y = 16'b1000000000010100;
        173: y = 16'b1000000000000010;
        174: y = 16'b1000000000001000;
        175: y = 16'b1000000000100110;
        176: y = 16'b1000000001011101;
        177: y = 16'b1000000010101011;
        178: y = 16'b1000000100010010;
        179: y = 16'b1000000110010001;
        180: y = 16'b1000001000101000;
        181: y = 16'b1000001011010110;
        182: y = 16'b1000001110011101;
        183: y = 16'b1000010001111011;
        184: y = 16'b1000010101110000;
        185: y = 16'b1000011001111100;
        186: y = 16'b1000011110100000;
        187: y = 16'b1000100011011010;
        188: y = 16'b1000101000101011;
        189: y = 16'b1000101110010010;
        190: y = 16'b1000110100001111;
        191: y = 16'b1000111010100010;
        192: y = 16'b1001000001001011;
        193: y = 16'b1001001000001000;
        194: y = 16'b1001001111011011;
        195: y = 16'b1001010111000010;
        196: y = 16'b1001011110111101;
        197: y = 16'b1001100111001100;
        198: y = 16'b1001101111101110;
        199: y = 16'b1001111000100011;
        200: y = 16'b1010000001101010;
        201: y = 16'b1010001011000100;
        202: y = 16'b1010010100110000;
        203: y = 16'b1010011110101100;
        204: y = 16'b1010101000111010;
        205: y = 16'b1010110011010111;
        206: y = 16'b1010111110000100;
        207: y = 16'b1011001001000001;
        208: y = 16'b1011010100001100;
        209: y = 16'b1011011111100110;
        210: y = 16'b1011101011001101;
        211: y = 16'b1011110111000001;
        212: y = 16'b1100000011000010;
        213: y = 16'b1100001111001111;
        214: y = 16'b1100011011100111;
        215: y = 16'b1100101000001010;
        216: y = 16'b1100110100110111;
        217: y = 16'b1101000001101110;
        218: y = 16'b1101001110101110;
        219: y = 16'b1101011011110110;
        220: y = 16'b1101101001000110;
        221: y = 16'b1101110110011101;
        222: y = 16'b1110000011111011;
        223: y = 16'b1110010001011110;
        224: y = 16'b1110011111000111;
        225: y = 16'b1110101100110100;
        226: y = 16'b1110111010100101;
        227: y = 16'b1111001000011010;
        228: y = 16'b1111010110010001;
        229: y = 16'b1111100100001010;
        230: y = 16'b1111110010000101;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=440.0Hz, Fs=96000Hz, 16-bit

module lut_A
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 217;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001110110000;
        2: y = 16'b0000011101100000;
        3: y = 16'b0000101100001110;
        4: y = 16'b0000111010111001;
        5: y = 16'b0001001001100010;
        6: y = 16'b0001011000000110;
        7: y = 16'b0001100110100110;
        8: y = 16'b0001110101000001;
        9: y = 16'b0010000011010101;
        10: y = 16'b0010010001100010;
        11: y = 16'b0010011111100111;
        12: y = 16'b0010101101100100;
        13: y = 16'b0010111011011000;
        14: y = 16'b0011001001000010;
        15: y = 16'b0011010110100001;
        16: y = 16'b0011100011110101;
        17: y = 16'b0011110000111100;
        18: y = 16'b0011111101110111;
        19: y = 16'b0100001010100100;
        20: y = 16'b0100010111000011;
        21: y = 16'b0100100011010100;
        22: y = 16'b0100101111010100;
        23: y = 16'b0100111011000101;
        24: y = 16'b0101000110100101;
        25: y = 16'b0101010001110100;
        26: y = 16'b0101011100110000;
        27: y = 16'b0101100111011010;
        28: y = 16'b0101110001110001;
        29: y = 16'b0101111011110100;
        30: y = 16'b0110000101100100;
        31: y = 16'b0110001110111110;
        32: y = 16'b0110011000000011;
        33: y = 16'b0110100000110011;
        34: y = 16'b0110101001001100;
        35: y = 16'b0110110001001111;
        36: y = 16'b0110111000111010;
        37: y = 16'b0111000000001111;
        38: y = 16'b0111000111001011;
        39: y = 16'b0111001101101111;
        40: y = 16'b0111010011111011;
        41: y = 16'b0111011001101110;
        42: y = 16'b0111011111000111;
        43: y = 16'b0111100100001000;
        44: y = 16'b0111101000101110;
        45: y = 16'b0111101100111010;
        46: y = 16'b0111110000101101;
        47: y = 16'b0111110100000100;
        48: y = 16'b0111110111000010;
        49: y = 16'b0111111001100100;
        50: y = 16'b0111111011101100;
        51: y = 16'b0111111101011000;
        52: y = 16'b0111111110101010;
        53: y = 16'b0111111111100000;
        54: y = 16'b0111111111111100;
        55: y = 16'b0111111111111100;
        56: y = 16'b0111111111100000;
        57: y = 16'b0111111110101010;
        58: y = 16'b0111111101011000;
        59: y = 16'b0111111011101100;
        60: y = 16'b0111111001100100;
        61: y = 16'b0111110111000010;
        62: y = 16'b0111110100000100;
        63: y = 16'b0111110000101101;
        64: y = 16'b0111101100111010;
        65: y = 16'b0111101000101110;
        66: y = 16'b0111100100001000;
        67: y = 16'b0111011111000111;
        68: y = 16'b0111011001101110;
        69: y = 16'b0111010011111011;
        70: y = 16'b0111001101101111;
        71: y = 16'b0111000111001011;
        72: y = 16'b0111000000001111;
        73: y = 16'b0110111000111010;
        74: y = 16'b0110110001001111;
        75: y = 16'b0110101001001100;
        76: y = 16'b0110100000110011;
        77: y = 16'b0110011000000011;
        78: y = 16'b0110001110111110;
        79: y = 16'b0110000101100100;
        80: y = 16'b0101111011110100;
        81: y = 16'b0101110001110001;
        82: y = 16'b0101100111011010;
        83: y = 16'b0101011100110000;
        84: y = 16'b0101010001110100;
        85: y = 16'b0101000110100101;
        86: y = 16'b0100111011000101;
        87: y = 16'b0100101111010100;
        88: y = 16'b0100100011010100;
        89: y = 16'b0100010111000011;
        90: y = 16'b0100001010100100;
        91: y = 16'b0011111101110111;
        92: y = 16'b0011110000111100;
        93: y = 16'b0011100011110101;
        94: y = 16'b0011010110100001;
        95: y = 16'b0011001001000010;
        96: y = 16'b0010111011011000;
        97: y = 16'b0010101101100100;
        98: y = 16'b0010011111100111;
        99: y = 16'b0010010001100010;
        100: y = 16'b0010000011010101;
        101: y = 16'b0001110101000001;
        102: y = 16'b0001100110100110;
        103: y = 16'b0001011000000110;
        104: y = 16'b0001001001100010;
        105: y = 16'b0000111010111001;
        106: y = 16'b0000101100001110;
        107: y = 16'b0000011101100000;
        108: y = 16'b0000001110110000;
        109: y = 16'b0000000000000000;
        110: y = 16'b1111110001010000;
        111: y = 16'b1111100010100000;
        112: y = 16'b1111010011110010;
        113: y = 16'b1111000101000111;
        114: y = 16'b1110110110011110;
        115: y = 16'b1110100111111010;
        116: y = 16'b1110011001011010;
        117: y = 16'b1110001010111111;
        118: y = 16'b1101111100101011;
        119: y = 16'b1101101110011110;
        120: y = 16'b1101100000011001;
        121: y = 16'b1101010010011100;
        122: y = 16'b1101000100101000;
        123: y = 16'b1100110110111110;
        124: y = 16'b1100101001011111;
        125: y = 16'b1100011100001011;
        126: y = 16'b1100001111000100;
        127: y = 16'b1100000010001001;
        128: y = 16'b1011110101011100;
        129: y = 16'b1011101000111101;
        130: y = 16'b1011011100101100;
        131: y = 16'b1011010000101100;
        132: y = 16'b1011000100111011;
        133: y = 16'b1010111001011011;
        134: y = 16'b1010101110001100;
        135: y = 16'b1010100011010000;
        136: y = 16'b1010011000100110;
        137: y = 16'b1010001110001111;
        138: y = 16'b1010000100001100;
        139: y = 16'b1001111010011100;
        140: y = 16'b1001110001000010;
        141: y = 16'b1001100111111101;
        142: y = 16'b1001011111001101;
        143: y = 16'b1001010110110100;
        144: y = 16'b1001001110110001;
        145: y = 16'b1001000111000110;
        146: y = 16'b1000111111110001;
        147: y = 16'b1000111000110101;
        148: y = 16'b1000110010010001;
        149: y = 16'b1000101100000101;
        150: y = 16'b1000100110010010;
        151: y = 16'b1000100000111001;
        152: y = 16'b1000011011111000;
        153: y = 16'b1000010111010010;
        154: y = 16'b1000010011000110;
        155: y = 16'b1000001111010011;
        156: y = 16'b1000001011111100;
        157: y = 16'b1000001000111110;
        158: y = 16'b1000000110011100;
        159: y = 16'b1000000100010100;
        160: y = 16'b1000000010101000;
        161: y = 16'b1000000001010110;
        162: y = 16'b1000000000100000;
        163: y = 16'b1000000000000100;
        164: y = 16'b1000000000000100;
        165: y = 16'b1000000000100000;
        166: y = 16'b1000000001010110;
        167: y = 16'b1000000010101000;
        168: y = 16'b1000000100010100;
        169: y = 16'b1000000110011100;
        170: y = 16'b1000001000111110;
        171: y = 16'b1000001011111100;
        172: y = 16'b1000001111010011;
        173: y = 16'b1000010011000110;
        174: y = 16'b1000010111010010;
        175: y = 16'b1000011011111000;
        176: y = 16'b1000100000111001;
        177: y = 16'b1000100110010010;
        178: y = 16'b1000101100000101;
        179: y = 16'b1000110010010001;
        180: y = 16'b1000111000110101;
        181: y = 16'b1000111111110001;
        182: y = 16'b1001000111000110;
        183: y = 16'b1001001110110001;
        184: y = 16'b1001010110110100;
        185: y = 16'b1001011111001101;
        186: y = 16'b1001100111111101;
        187: y = 16'b1001110001000010;
        188: y = 16'b1001111010011100;
        189: y = 16'b1010000100001100;
        190: y = 16'b1010001110001111;
        191: y = 16'b1010011000100110;
        192: y = 16'b1010100011010000;
        193: y = 16'b1010101110001100;
        194: y = 16'b1010111001011011;
        195: y = 16'b1011000100111011;
        196: y = 16'b1011010000101100;
        197: y = 16'b1011011100101100;
        198: y = 16'b1011101000111101;
        199: y = 16'b1011110101011100;
        200: y = 16'b1100000010001001;
        201: y = 16'b1100001111000100;
        202: y = 16'b1100011100001011;
        203: y = 16'b1100101001011111;
        204: y = 16'b1100110110111110;
        205: y = 16'b1101000100101000;
        206: y = 16'b1101010010011100;
        207: y = 16'b1101100000011001;
        208: y = 16'b1101101110011110;
        209: y = 16'b1101111100101011;
        210: y = 16'b1110001010111111;
        211: y = 16'b1110011001011010;
        212: y = 16'b1110100111111010;
        213: y = 16'b1110110110011110;
        214: y = 16'b1111000101000111;
        215: y = 16'b1111010011110010;
        216: y = 16'b1111100010100000;
        217: y = 16'b1111110001010000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=466.16Hz, Fs=96000Hz, 16-bit

module lut_As
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 204;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001111101100;
        2: y = 16'b0000011111010111;
        3: y = 16'b0000101111000001;
        4: y = 16'b0000111110100111;
        5: y = 16'b0001001110001010;
        6: y = 16'b0001011101101000;
        7: y = 16'b0001101101000000;
        8: y = 16'b0001111100010010;
        9: y = 16'b0010001011011100;
        10: y = 16'b0010011010011110;
        11: y = 16'b0010101001010111;
        12: y = 16'b0010111000000110;
        13: y = 16'b0011000110101001;
        14: y = 16'b0011010101000001;
        15: y = 16'b0011100011001011;
        16: y = 16'b0011110001001000;
        17: y = 16'b0011111110110111;
        18: y = 16'b0100001100010110;
        19: y = 16'b0100011001100101;
        20: y = 16'b0100100110100011;
        21: y = 16'b0100110011010000;
        22: y = 16'b0100111111101010;
        23: y = 16'b0101001011110001;
        24: y = 16'b0101010111100100;
        25: y = 16'b0101100011000010;
        26: y = 16'b0101101110001011;
        27: y = 16'b0101111000111101;
        28: y = 16'b0110000011011010;
        29: y = 16'b0110001101011110;
        30: y = 16'b0110010111001011;
        31: y = 16'b0110100000100000;
        32: y = 16'b0110101001011011;
        33: y = 16'b0110110001111101;
        34: y = 16'b0110111010000101;
        35: y = 16'b0111000001110010;
        36: y = 16'b0111001001000100;
        37: y = 16'b0111001111111011;
        38: y = 16'b0111010110010110;
        39: y = 16'b0111011100010100;
        40: y = 16'b0111100001110110;
        41: y = 16'b0111100110111011;
        42: y = 16'b0111101011100011;
        43: y = 16'b0111101111101101;
        44: y = 16'b0111110011011001;
        45: y = 16'b0111110110101000;
        46: y = 16'b0111111001011000;
        47: y = 16'b0111111011101001;
        48: y = 16'b0111111101011101;
        49: y = 16'b0111111110110001;
        50: y = 16'b0111111111100111;
        51: y = 16'b0111111111111110;
        52: y = 16'b0111111111110110;
        53: y = 16'b0111111111010000;
        54: y = 16'b0111111110001011;
        55: y = 16'b0111111100100111;
        56: y = 16'b0111111010100100;
        57: y = 16'b0111111000000011;
        58: y = 16'b0111110101000100;
        59: y = 16'b0111110001100111;
        60: y = 16'b0111101101101100;
        61: y = 16'b0111101001010011;
        62: y = 16'b0111100100011100;
        63: y = 16'b0111011111001001;
        64: y = 16'b0111011001011001;
        65: y = 16'b0111010011001100;
        66: y = 16'b0111001100100011;
        67: y = 16'b0111000101011111;
        68: y = 16'b0110111101111111;
        69: y = 16'b0110110110000100;
        70: y = 16'b0110101101101111;
        71: y = 16'b0110100101000001;
        72: y = 16'b0110011011111001;
        73: y = 16'b0110010010011000;
        74: y = 16'b0110001000011111;
        75: y = 16'b0101111110001110;
        76: y = 16'b0101110011100111;
        77: y = 16'b0101101000101001;
        78: y = 16'b0101011101010101;
        79: y = 16'b0101010001101101;
        80: y = 16'b0101000101110000;
        81: y = 16'b0100111001011111;
        82: y = 16'b0100101100111100;
        83: y = 16'b0100100000000111;
        84: y = 16'b0100010011000000;
        85: y = 16'b0100000101101001;
        86: y = 16'b0011111000000010;
        87: y = 16'b0011101010001100;
        88: y = 16'b0011011100001000;
        89: y = 16'b0011001101110110;
        90: y = 16'b0010111111011001;
        91: y = 16'b0010110000110000;
        92: y = 16'b0010100001111100;
        93: y = 16'b0010010010111111;
        94: y = 16'b0010000011111000;
        95: y = 16'b0001110100101010;
        96: y = 16'b0001100101010101;
        97: y = 16'b0001010101111010;
        98: y = 16'b0001000110011001;
        99: y = 16'b0000110110110100;
        100: y = 16'b0000100111001100;
        101: y = 16'b0000010111100010;
        102: y = 16'b0000000111110110;
        103: y = 16'b1111111000001010;
        104: y = 16'b1111101000011110;
        105: y = 16'b1111011000110100;
        106: y = 16'b1111001001001100;
        107: y = 16'b1110111001100111;
        108: y = 16'b1110101010000110;
        109: y = 16'b1110011010101011;
        110: y = 16'b1110001011010110;
        111: y = 16'b1101111100001000;
        112: y = 16'b1101101101000001;
        113: y = 16'b1101011110000100;
        114: y = 16'b1101001111010000;
        115: y = 16'b1101000000100111;
        116: y = 16'b1100110010001010;
        117: y = 16'b1100100011111000;
        118: y = 16'b1100010101110100;
        119: y = 16'b1100000111111110;
        120: y = 16'b1011111010010111;
        121: y = 16'b1011101101000000;
        122: y = 16'b1011011111111001;
        123: y = 16'b1011010011000100;
        124: y = 16'b1011000110100001;
        125: y = 16'b1010111010010000;
        126: y = 16'b1010101110010011;
        127: y = 16'b1010100010101011;
        128: y = 16'b1010010111010111;
        129: y = 16'b1010001100011001;
        130: y = 16'b1010000001110010;
        131: y = 16'b1001110111100001;
        132: y = 16'b1001101101101000;
        133: y = 16'b1001100100000111;
        134: y = 16'b1001011010111111;
        135: y = 16'b1001010010010001;
        136: y = 16'b1001001001111100;
        137: y = 16'b1001000010000001;
        138: y = 16'b1000111010100001;
        139: y = 16'b1000110011011101;
        140: y = 16'b1000101100110100;
        141: y = 16'b1000100110100111;
        142: y = 16'b1000100000110111;
        143: y = 16'b1000011011100100;
        144: y = 16'b1000010110101101;
        145: y = 16'b1000010010010100;
        146: y = 16'b1000001110011001;
        147: y = 16'b1000001010111100;
        148: y = 16'b1000000111111101;
        149: y = 16'b1000000101011100;
        150: y = 16'b1000000011011001;
        151: y = 16'b1000000001110101;
        152: y = 16'b1000000000110000;
        153: y = 16'b1000000000001010;
        154: y = 16'b1000000000000010;
        155: y = 16'b1000000000011001;
        156: y = 16'b1000000001001111;
        157: y = 16'b1000000010100011;
        158: y = 16'b1000000100010111;
        159: y = 16'b1000000110101000;
        160: y = 16'b1000001001011000;
        161: y = 16'b1000001100100111;
        162: y = 16'b1000010000010011;
        163: y = 16'b1000010100011101;
        164: y = 16'b1000011001000101;
        165: y = 16'b1000011110001010;
        166: y = 16'b1000100011101100;
        167: y = 16'b1000101001101010;
        168: y = 16'b1000110000000101;
        169: y = 16'b1000110110111100;
        170: y = 16'b1000111110001110;
        171: y = 16'b1001000101111011;
        172: y = 16'b1001001110000011;
        173: y = 16'b1001010110100101;
        174: y = 16'b1001011111100000;
        175: y = 16'b1001101000110101;
        176: y = 16'b1001110010100010;
        177: y = 16'b1001111100100110;
        178: y = 16'b1010000111000011;
        179: y = 16'b1010010001110101;
        180: y = 16'b1010011100111110;
        181: y = 16'b1010101000011100;
        182: y = 16'b1010110100001111;
        183: y = 16'b1011000000010110;
        184: y = 16'b1011001100110000;
        185: y = 16'b1011011001011101;
        186: y = 16'b1011100110011011;
        187: y = 16'b1011110011101010;
        188: y = 16'b1100000001001001;
        189: y = 16'b1100001110111000;
        190: y = 16'b1100011100110101;
        191: y = 16'b1100101010111111;
        192: y = 16'b1100111001010111;
        193: y = 16'b1101000111111010;
        194: y = 16'b1101010110101001;
        195: y = 16'b1101100101100010;
        196: y = 16'b1101110100100100;
        197: y = 16'b1110000011101110;
        198: y = 16'b1110010011000000;
        199: y = 16'b1110100010011000;
        200: y = 16'b1110110001110110;
        201: y = 16'b1111000001011001;
        202: y = 16'b1111010000111111;
        203: y = 16'b1111100000101001;
        204: y = 16'b1111110000010100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=493.88Hz, Fs=96000Hz, 16-bit

module lut_B
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 193;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000010000100101;
        2: y = 16'b0000100001001001;
        3: y = 16'b0000110001101011;
        4: y = 16'b0001000010001001;
        5: y = 16'b0001010010100011;
        6: y = 16'b0001100010110111;
        7: y = 16'b0001110011000101;
        8: y = 16'b0010000011001011;
        9: y = 16'b0010010011001001;
        10: y = 16'b0010100010111100;
        11: y = 16'b0010110010100100;
        12: y = 16'b0011000010000001;
        13: y = 16'b0011010001010000;
        14: y = 16'b0011100000010010;
        15: y = 16'b0011101111000100;
        16: y = 16'b0011111101100110;
        17: y = 16'b0100001011110111;
        18: y = 16'b0100011001110111;
        19: y = 16'b0100100111100011;
        20: y = 16'b0100110100111011;
        21: y = 16'b0101000001111111;
        22: y = 16'b0101001110101101;
        23: y = 16'b0101011011000101;
        24: y = 16'b0101100111000101;
        25: y = 16'b0101110010101110;
        26: y = 16'b0101111101111101;
        27: y = 16'b0110001000110011;
        28: y = 16'b0110010011001110;
        29: y = 16'b0110011101001111;
        30: y = 16'b0110100110110011;
        31: y = 16'b0110101111111011;
        32: y = 16'b0110111000100111;
        33: y = 16'b0111000000110100;
        34: y = 16'b0111001000100100;
        35: y = 16'b0111001111110101;
        36: y = 16'b0111010110100110;
        37: y = 16'b0111011100111000;
        38: y = 16'b0111100010101010;
        39: y = 16'b0111100111111100;
        40: y = 16'b0111101100101101;
        41: y = 16'b0111110000111101;
        42: y = 16'b0111110100101100;
        43: y = 16'b0111110111111001;
        44: y = 16'b0111111010100100;
        45: y = 16'b0111111100101101;
        46: y = 16'b0111111110010100;
        47: y = 16'b0111111111011000;
        48: y = 16'b0111111111111011;
        49: y = 16'b0111111111111011;
        50: y = 16'b0111111111011000;
        51: y = 16'b0111111110010100;
        52: y = 16'b0111111100101101;
        53: y = 16'b0111111010100100;
        54: y = 16'b0111110111111001;
        55: y = 16'b0111110100101100;
        56: y = 16'b0111110000111101;
        57: y = 16'b0111101100101101;
        58: y = 16'b0111100111111100;
        59: y = 16'b0111100010101010;
        60: y = 16'b0111011100111000;
        61: y = 16'b0111010110100110;
        62: y = 16'b0111001111110101;
        63: y = 16'b0111001000100100;
        64: y = 16'b0111000000110100;
        65: y = 16'b0110111000100111;
        66: y = 16'b0110101111111011;
        67: y = 16'b0110100110110011;
        68: y = 16'b0110011101001111;
        69: y = 16'b0110010011001110;
        70: y = 16'b0110001000110011;
        71: y = 16'b0101111101111101;
        72: y = 16'b0101110010101110;
        73: y = 16'b0101100111000101;
        74: y = 16'b0101011011000101;
        75: y = 16'b0101001110101101;
        76: y = 16'b0101000001111111;
        77: y = 16'b0100110100111011;
        78: y = 16'b0100100111100011;
        79: y = 16'b0100011001110111;
        80: y = 16'b0100001011110111;
        81: y = 16'b0011111101100110;
        82: y = 16'b0011101111000100;
        83: y = 16'b0011100000010010;
        84: y = 16'b0011010001010000;
        85: y = 16'b0011000010000001;
        86: y = 16'b0010110010100100;
        87: y = 16'b0010100010111100;
        88: y = 16'b0010010011001001;
        89: y = 16'b0010000011001011;
        90: y = 16'b0001110011000101;
        91: y = 16'b0001100010110111;
        92: y = 16'b0001010010100011;
        93: y = 16'b0001000010001001;
        94: y = 16'b0000110001101011;
        95: y = 16'b0000100001001001;
        96: y = 16'b0000010000100101;
        97: y = 16'b0000000000000000;
        98: y = 16'b1111101111011011;
        99: y = 16'b1111011110110111;
        100: y = 16'b1111001110010101;
        101: y = 16'b1110111101110111;
        102: y = 16'b1110101101011101;
        103: y = 16'b1110011101001001;
        104: y = 16'b1110001100111011;
        105: y = 16'b1101111100110101;
        106: y = 16'b1101101100110111;
        107: y = 16'b1101011101000100;
        108: y = 16'b1101001101011100;
        109: y = 16'b1100111101111111;
        110: y = 16'b1100101110110000;
        111: y = 16'b1100011111101110;
        112: y = 16'b1100010000111100;
        113: y = 16'b1100000010011010;
        114: y = 16'b1011110100001001;
        115: y = 16'b1011100110001001;
        116: y = 16'b1011011000011101;
        117: y = 16'b1011001011000101;
        118: y = 16'b1010111110000001;
        119: y = 16'b1010110001010011;
        120: y = 16'b1010100100111011;
        121: y = 16'b1010011000111011;
        122: y = 16'b1010001101010010;
        123: y = 16'b1010000010000011;
        124: y = 16'b1001110111001101;
        125: y = 16'b1001101100110010;
        126: y = 16'b1001100010110001;
        127: y = 16'b1001011001001101;
        128: y = 16'b1001010000000101;
        129: y = 16'b1001000111011001;
        130: y = 16'b1000111111001100;
        131: y = 16'b1000110111011100;
        132: y = 16'b1000110000001011;
        133: y = 16'b1000101001011010;
        134: y = 16'b1000100011001000;
        135: y = 16'b1000011101010110;
        136: y = 16'b1000011000000100;
        137: y = 16'b1000010011010011;
        138: y = 16'b1000001111000011;
        139: y = 16'b1000001011010100;
        140: y = 16'b1000001000000111;
        141: y = 16'b1000000101011100;
        142: y = 16'b1000000011010011;
        143: y = 16'b1000000001101100;
        144: y = 16'b1000000000101000;
        145: y = 16'b1000000000000101;
        146: y = 16'b1000000000000101;
        147: y = 16'b1000000000101000;
        148: y = 16'b1000000001101100;
        149: y = 16'b1000000011010011;
        150: y = 16'b1000000101011100;
        151: y = 16'b1000001000000111;
        152: y = 16'b1000001011010100;
        153: y = 16'b1000001111000011;
        154: y = 16'b1000010011010011;
        155: y = 16'b1000011000000100;
        156: y = 16'b1000011101010110;
        157: y = 16'b1000100011001000;
        158: y = 16'b1000101001011010;
        159: y = 16'b1000110000001011;
        160: y = 16'b1000110111011100;
        161: y = 16'b1000111111001100;
        162: y = 16'b1001000111011001;
        163: y = 16'b1001010000000101;
        164: y = 16'b1001011001001101;
        165: y = 16'b1001100010110001;
        166: y = 16'b1001101100110010;
        167: y = 16'b1001110111001101;
        168: y = 16'b1010000010000011;
        169: y = 16'b1010001101010010;
        170: y = 16'b1010011000111011;
        171: y = 16'b1010100100111011;
        172: y = 16'b1010110001010011;
        173: y = 16'b1010111110000001;
        174: y = 16'b1011001011000101;
        175: y = 16'b1011011000011101;
        176: y = 16'b1011100110001001;
        177: y = 16'b1011110100001001;
        178: y = 16'b1100000010011010;
        179: y = 16'b1100010000111100;
        180: y = 16'b1100011111101110;
        181: y = 16'b1100101110110000;
        182: y = 16'b1100111101111111;
        183: y = 16'b1101001101011100;
        184: y = 16'b1101011101000100;
        185: y = 16'b1101101100110111;
        186: y = 16'b1101111100110101;
        187: y = 16'b1110001100111011;
        188: y = 16'b1110011101001001;
        189: y = 16'b1110101101011101;
        190: y = 16'b1110111101110111;
        191: y = 16'b1111001110010101;
        192: y = 16'b1111011110110111;
        193: y = 16'b1111101111011011;
        default: y = 16'b0;
        endcase

endmodule

