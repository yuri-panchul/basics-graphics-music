`include "config.svh"

module lab_top
# (
    parameter  clk_mhz       = 50,
               w_key         = 4,
               w_sw          = 8,
               w_led         = 8,
               w_digit       = 8,
               w_gpio        = 100,

               screen_width  = 640,
               screen_height = 480,

               w_red         = 4,
               w_green       = 4,
               w_blue        = 4,

               w_x           = $clog2 ( screen_width  ),
               w_y           = $clog2 ( screen_height )
)
(
    input                        clk,
    input                        slow_clk,
    input                        rst,

    // Keys, switches, LEDs

    input        [w_key   - 1:0] key,
    input        [w_sw    - 1:0] sw,
    output logic [w_led   - 1:0] led,

    // A dynamic seven-segment display

    output logic [          7:0] abcdefgh,
    output logic [w_digit - 1:0] digit,

    // Graphics

    input        [w_x     - 1:0] x,
    input        [w_y     - 1:0] y,

    output logic [w_red   - 1:0] red,
    output logic [w_green - 1:0] green,
    output logic [w_blue  - 1:0] blue,

    // Microphone, sound output and UART

    input        [         23:0] mic,
    output       [         15:0] sound,

    input                        uart_rx,
    output                       uart_tx,

    // General-purpose Input/Output

    inout        [w_gpio  - 1:0] gpio
);

    //------------------------------------------------------------------------

       assign led        = '0;
       assign abcdefgh   = '0;
       assign digit      = '0;
    // assign red        = '0;
    // assign green      = '0;
    // assign blue       = '0;
       assign sound      = '0;
       assign uart_tx    = '1;

    //------------------------------------------------------------------------
    //
    //  NOTE! Since Maker Faire examples are for absolute beginners,
    //  we are using simplified, more relaxed Verilog style.
    //  For example, "100" instead of "w_x' (100)" or  "screen_width / 2".
    //
    //------------------------------------------------------------------------

    logic [9:0] w;

    always_comb
    begin
        red   = 0;
        green = 0;
        blue  = 0;

        if (x > 100 & y > 100 & x < 150 & y < 200)
        begin
            red   = key [0] ? 30 : 0;
            green = key [1] ? 30 : 0;
            blue  = key [2] ? 30 : 0;
        end

        if (key [4])
            w = 200;
        else
            w = 50;

        if (x > 200 & y > 0 & x < 200 + w & y < 100)
            green = 30;
    end

endmodule
