// y(t) = sin(2*pi*F*t), F=261.63Hz, Fs=64453Hz, 16-bit

module lut_C
(
    input        [ 7:0] x,
    output       [ 7:0] x_max,
    output logic [15:0] y
);

    assign x_max = 245;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000000110100010;
        2: y = 16'b0000001101000101;
        3: y = 16'b0000010011100110;
        4: y = 16'b0000011010000111;
        5: y = 16'b0000100000100111;
        6: y = 16'b0000100111000101;
        7: y = 16'b0000101101100010;
        8: y = 16'b0000110011111100;
        9: y = 16'b0000111010010101;
        10: y = 16'b0001000000101011;
        11: y = 16'b0001000110111111;
        12: y = 16'b0001001101001111;
        13: y = 16'b0001010011011100;
        14: y = 16'b0001011001100110;
        15: y = 16'b0001011111101100;
        16: y = 16'b0001100101101110;
        17: y = 16'b0001101011101100;
        18: y = 16'b0001110001100101;
        19: y = 16'b0001110111011010;
        20: y = 16'b0001111101001010;
        21: y = 16'b0010000010110100;
        22: y = 16'b0010001000011001;
        23: y = 16'b0010001101111000;
        24: y = 16'b0010010011010001;
        25: y = 16'b0010011000100101;
        26: y = 16'b0010011101110001;
        27: y = 16'b0010100010111000;
        28: y = 16'b0010100111110111;
        29: y = 16'b0010101100101111;
        30: y = 16'b0010110001100001;
        31: y = 16'b0010110110001010;
        32: y = 16'b0010111010101100;
        33: y = 16'b0010111111000111;
        34: y = 16'b0011000011011001;
        35: y = 16'b0011000111100011;
        36: y = 16'b0011001011100101;
        37: y = 16'b0011001111011111;
        38: y = 16'b0011010011001111;
        39: y = 16'b0011010110110111;
        40: y = 16'b0011011010010110;
        41: y = 16'b0011011101101100;
        42: y = 16'b0011100000111001;
        43: y = 16'b0011100011111100;
        44: y = 16'b0011100110110110;
        45: y = 16'b0011101001100110;
        46: y = 16'b0011101100001100;
        47: y = 16'b0011101110101000;
        48: y = 16'b0011110000111011;
        49: y = 16'b0011110011000011;
        50: y = 16'b0011110101000001;
        51: y = 16'b0011110110110101;
        52: y = 16'b0011111000011111;
        53: y = 16'b0011111001111110;
        54: y = 16'b0011111011010011;
        55: y = 16'b0011111100011110;
        56: y = 16'b0011111101011110;
        57: y = 16'b0011111110010011;
        58: y = 16'b0011111110111110;
        59: y = 16'b0011111111011110;
        60: y = 16'b0011111111110011;
        61: y = 16'b0011111111111110;
        62: y = 16'b0011111111111110;
        63: y = 16'b0011111111110011;
        64: y = 16'b0011111111011110;
        65: y = 16'b0011111110111110;
        66: y = 16'b0011111110010011;
        67: y = 16'b0011111101011110;
        68: y = 16'b0011111100011110;
        69: y = 16'b0011111011010011;
        70: y = 16'b0011111001111110;
        71: y = 16'b0011111000011111;
        72: y = 16'b0011110110110101;
        73: y = 16'b0011110101000001;
        74: y = 16'b0011110011000011;
        75: y = 16'b0011110000111011;
        76: y = 16'b0011101110101000;
        77: y = 16'b0011101100001100;
        78: y = 16'b0011101001100110;
        79: y = 16'b0011100110110110;
        80: y = 16'b0011100011111100;
        81: y = 16'b0011100000111001;
        82: y = 16'b0011011101101100;
        83: y = 16'b0011011010010110;
        84: y = 16'b0011010110110111;
        85: y = 16'b0011010011001111;
        86: y = 16'b0011001111011111;
        87: y = 16'b0011001011100101;
        88: y = 16'b0011000111100011;
        89: y = 16'b0011000011011001;
        90: y = 16'b0010111111000111;
        91: y = 16'b0010111010101100;
        92: y = 16'b0010110110001010;
        93: y = 16'b0010110001100001;
        94: y = 16'b0010101100101111;
        95: y = 16'b0010100111110111;
        96: y = 16'b0010100010111000;
        97: y = 16'b0010011101110001;
        98: y = 16'b0010011000100101;
        99: y = 16'b0010010011010001;
        100: y = 16'b0010001101111000;
        101: y = 16'b0010001000011001;
        102: y = 16'b0010000010110100;
        103: y = 16'b0001111101001010;
        104: y = 16'b0001110111011010;
        105: y = 16'b0001110001100101;
        106: y = 16'b0001101011101100;
        107: y = 16'b0001100101101110;
        108: y = 16'b0001011111101100;
        109: y = 16'b0001011001100110;
        110: y = 16'b0001010011011100;
        111: y = 16'b0001001101001111;
        112: y = 16'b0001000110111111;
        113: y = 16'b0001000000101011;
        114: y = 16'b0000111010010101;
        115: y = 16'b0000110011111100;
        116: y = 16'b0000101101100010;
        117: y = 16'b0000100111000101;
        118: y = 16'b0000100000100111;
        119: y = 16'b0000011010000111;
        120: y = 16'b0000010011100110;
        121: y = 16'b0000001101000101;
        122: y = 16'b0000000110100010;
        123: y = 16'b0000000000000000;
        124: y = 16'b1111111001011110;
        125: y = 16'b1111110010111011;
        126: y = 16'b1111101100011010;
        127: y = 16'b1111100101111001;
        128: y = 16'b1111011111011001;
        129: y = 16'b1111011000111011;
        130: y = 16'b1111010010011110;
        131: y = 16'b1111001100000100;
        132: y = 16'b1111000101101011;
        133: y = 16'b1110111111010101;
        134: y = 16'b1110111001000001;
        135: y = 16'b1110110010110001;
        136: y = 16'b1110101100100100;
        137: y = 16'b1110100110011010;
        138: y = 16'b1110100000010100;
        139: y = 16'b1110011010010010;
        140: y = 16'b1110010100010100;
        141: y = 16'b1110001110011011;
        142: y = 16'b1110001000100110;
        143: y = 16'b1110000010110110;
        144: y = 16'b1101111101001100;
        145: y = 16'b1101110111100111;
        146: y = 16'b1101110010001000;
        147: y = 16'b1101101100101111;
        148: y = 16'b1101100111011011;
        149: y = 16'b1101100010001111;
        150: y = 16'b1101011101001000;
        151: y = 16'b1101011000001001;
        152: y = 16'b1101010011010001;
        153: y = 16'b1101001110011111;
        154: y = 16'b1101001001110110;
        155: y = 16'b1101000101010100;
        156: y = 16'b1101000000111001;
        157: y = 16'b1100111100100111;
        158: y = 16'b1100111000011101;
        159: y = 16'b1100110100011011;
        160: y = 16'b1100110000100001;
        161: y = 16'b1100101100110001;
        162: y = 16'b1100101001001001;
        163: y = 16'b1100100101101010;
        164: y = 16'b1100100010010100;
        165: y = 16'b1100011111000111;
        166: y = 16'b1100011100000100;
        167: y = 16'b1100011001001010;
        168: y = 16'b1100010110011010;
        169: y = 16'b1100010011110100;
        170: y = 16'b1100010001011000;
        171: y = 16'b1100001111000101;
        172: y = 16'b1100001100111101;
        173: y = 16'b1100001010111111;
        174: y = 16'b1100001001001011;
        175: y = 16'b1100000111100001;
        176: y = 16'b1100000110000010;
        177: y = 16'b1100000100101101;
        178: y = 16'b1100000011100010;
        179: y = 16'b1100000010100010;
        180: y = 16'b1100000001101101;
        181: y = 16'b1100000001000010;
        182: y = 16'b1100000000100010;
        183: y = 16'b1100000000001101;
        184: y = 16'b1100000000000010;
        185: y = 16'b1100000000000010;
        186: y = 16'b1100000000001101;
        187: y = 16'b1100000000100010;
        188: y = 16'b1100000001000010;
        189: y = 16'b1100000001101101;
        190: y = 16'b1100000010100010;
        191: y = 16'b1100000011100010;
        192: y = 16'b1100000100101101;
        193: y = 16'b1100000110000010;
        194: y = 16'b1100000111100001;
        195: y = 16'b1100001001001011;
        196: y = 16'b1100001010111111;
        197: y = 16'b1100001100111101;
        198: y = 16'b1100001111000101;
        199: y = 16'b1100010001011000;
        200: y = 16'b1100010011110100;
        201: y = 16'b1100010110011010;
        202: y = 16'b1100011001001010;
        203: y = 16'b1100011100000100;
        204: y = 16'b1100011111000111;
        205: y = 16'b1100100010010100;
        206: y = 16'b1100100101101010;
        207: y = 16'b1100101001001001;
        208: y = 16'b1100101100110001;
        209: y = 16'b1100110000100001;
        210: y = 16'b1100110100011011;
        211: y = 16'b1100111000011101;
        212: y = 16'b1100111100100111;
        213: y = 16'b1101000000111001;
        214: y = 16'b1101000101010100;
        215: y = 16'b1101001001110110;
        216: y = 16'b1101001110011111;
        217: y = 16'b1101010011010001;
        218: y = 16'b1101011000001001;
        219: y = 16'b1101011101001000;
        220: y = 16'b1101100010001111;
        221: y = 16'b1101100111011011;
        222: y = 16'b1101101100101111;
        223: y = 16'b1101110010001000;
        224: y = 16'b1101110111100111;
        225: y = 16'b1101111101001100;
        226: y = 16'b1110000010110110;
        227: y = 16'b1110001000100110;
        228: y = 16'b1110001110011011;
        229: y = 16'b1110010100010100;
        230: y = 16'b1110011010010010;
        231: y = 16'b1110100000010100;
        232: y = 16'b1110100110011010;
        233: y = 16'b1110101100100100;
        234: y = 16'b1110110010110001;
        235: y = 16'b1110111001000001;
        236: y = 16'b1110111111010101;
        237: y = 16'b1111000101101011;
        238: y = 16'b1111001100000100;
        239: y = 16'b1111010010011110;
        240: y = 16'b1111011000111011;
        241: y = 16'b1111011111011001;
        242: y = 16'b1111100101111001;
        243: y = 16'b1111101100011010;
        244: y = 16'b1111110010111011;
        245: y = 16'b1111111001011110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=277.18Hz, Fs=64453Hz, 16-bit

module lut_Cs
(
    input        [ 7:0] x,
    output       [ 7:0] x_max,
    output logic [15:0] y
);

    assign x_max = 231;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000000110111100;
        2: y = 16'b0000001101110111;
        3: y = 16'b0000010100110010;
        4: y = 16'b0000011011101011;
        5: y = 16'b0000100010100100;
        6: y = 16'b0000101001011010;
        7: y = 16'b0000110000001111;
        8: y = 16'b0000110111000010;
        9: y = 16'b0000111101110010;
        10: y = 16'b0001000100011111;
        11: y = 16'b0001001011001001;
        12: y = 16'b0001010001101111;
        13: y = 16'b0001011000010010;
        14: y = 16'b0001011110110000;
        15: y = 16'b0001100101001010;
        16: y = 16'b0001101011011111;
        17: y = 16'b0001110001101111;
        18: y = 16'b0001110111111010;
        19: y = 16'b0001111101111111;
        20: y = 16'b0010000011111110;
        21: y = 16'b0010001001110111;
        22: y = 16'b0010001111101010;
        23: y = 16'b0010010101010110;
        24: y = 16'b0010011010111011;
        25: y = 16'b0010100000011000;
        26: y = 16'b0010100101101110;
        27: y = 16'b0010101010111100;
        28: y = 16'b0010110000000011;
        29: y = 16'b0010110101000001;
        30: y = 16'b0010111001110110;
        31: y = 16'b0010111110100011;
        32: y = 16'b0011000011000111;
        33: y = 16'b0011000111100001;
        34: y = 16'b0011001011110010;
        35: y = 16'b0011001111111010;
        36: y = 16'b0011010011111000;
        37: y = 16'b0011010111101100;
        38: y = 16'b0011011011010110;
        39: y = 16'b0011011110110101;
        40: y = 16'b0011100010001011;
        41: y = 16'b0011100101010101;
        42: y = 16'b0011101000010101;
        43: y = 16'b0011101011001010;
        44: y = 16'b0011101101110011;
        45: y = 16'b0011110000010010;
        46: y = 16'b0011110010100101;
        47: y = 16'b0011110100101101;
        48: y = 16'b0011110110101010;
        49: y = 16'b0011111000011011;
        50: y = 16'b0011111010000000;
        51: y = 16'b0011111011011001;
        52: y = 16'b0011111100100111;
        53: y = 16'b0011111101101001;
        54: y = 16'b0011111110011111;
        55: y = 16'b0011111111001001;
        56: y = 16'b0011111111100111;
        57: y = 16'b0011111111111001;
        58: y = 16'b0011111111111111;
        59: y = 16'b0011111111111001;
        60: y = 16'b0011111111100111;
        61: y = 16'b0011111111001001;
        62: y = 16'b0011111110011111;
        63: y = 16'b0011111101101001;
        64: y = 16'b0011111100100111;
        65: y = 16'b0011111011011001;
        66: y = 16'b0011111010000000;
        67: y = 16'b0011111000011011;
        68: y = 16'b0011110110101010;
        69: y = 16'b0011110100101101;
        70: y = 16'b0011110010100101;
        71: y = 16'b0011110000010010;
        72: y = 16'b0011101101110011;
        73: y = 16'b0011101011001010;
        74: y = 16'b0011101000010101;
        75: y = 16'b0011100101010101;
        76: y = 16'b0011100010001011;
        77: y = 16'b0011011110110101;
        78: y = 16'b0011011011010110;
        79: y = 16'b0011010111101100;
        80: y = 16'b0011010011111000;
        81: y = 16'b0011001111111010;
        82: y = 16'b0011001011110010;
        83: y = 16'b0011000111100001;
        84: y = 16'b0011000011000111;
        85: y = 16'b0010111110100011;
        86: y = 16'b0010111001110110;
        87: y = 16'b0010110101000001;
        88: y = 16'b0010110000000011;
        89: y = 16'b0010101010111100;
        90: y = 16'b0010100101101110;
        91: y = 16'b0010100000011000;
        92: y = 16'b0010011010111011;
        93: y = 16'b0010010101010110;
        94: y = 16'b0010001111101010;
        95: y = 16'b0010001001110111;
        96: y = 16'b0010000011111110;
        97: y = 16'b0001111101111111;
        98: y = 16'b0001110111111010;
        99: y = 16'b0001110001101111;
        100: y = 16'b0001101011011111;
        101: y = 16'b0001100101001010;
        102: y = 16'b0001011110110000;
        103: y = 16'b0001011000010010;
        104: y = 16'b0001010001101111;
        105: y = 16'b0001001011001001;
        106: y = 16'b0001000100011111;
        107: y = 16'b0000111101110010;
        108: y = 16'b0000110111000010;
        109: y = 16'b0000110000001111;
        110: y = 16'b0000101001011010;
        111: y = 16'b0000100010100100;
        112: y = 16'b0000011011101011;
        113: y = 16'b0000010100110010;
        114: y = 16'b0000001101110111;
        115: y = 16'b0000000110111100;
        116: y = 16'b0000000000000000;
        117: y = 16'b1111111001000100;
        118: y = 16'b1111110010001001;
        119: y = 16'b1111101011001110;
        120: y = 16'b1111100100010101;
        121: y = 16'b1111011101011100;
        122: y = 16'b1111010110100110;
        123: y = 16'b1111001111110001;
        124: y = 16'b1111001000111110;
        125: y = 16'b1111000010001110;
        126: y = 16'b1110111011100001;
        127: y = 16'b1110110100110111;
        128: y = 16'b1110101110010001;
        129: y = 16'b1110100111101110;
        130: y = 16'b1110100001010000;
        131: y = 16'b1110011010110110;
        132: y = 16'b1110010100100001;
        133: y = 16'b1110001110010001;
        134: y = 16'b1110001000000110;
        135: y = 16'b1110000010000001;
        136: y = 16'b1101111100000010;
        137: y = 16'b1101110110001001;
        138: y = 16'b1101110000010110;
        139: y = 16'b1101101010101010;
        140: y = 16'b1101100101000101;
        141: y = 16'b1101011111101000;
        142: y = 16'b1101011010010010;
        143: y = 16'b1101010101000100;
        144: y = 16'b1101001111111101;
        145: y = 16'b1101001010111111;
        146: y = 16'b1101000110001010;
        147: y = 16'b1101000001011101;
        148: y = 16'b1100111100111001;
        149: y = 16'b1100111000011111;
        150: y = 16'b1100110100001110;
        151: y = 16'b1100110000000110;
        152: y = 16'b1100101100001000;
        153: y = 16'b1100101000010100;
        154: y = 16'b1100100100101010;
        155: y = 16'b1100100001001011;
        156: y = 16'b1100011101110101;
        157: y = 16'b1100011010101011;
        158: y = 16'b1100010111101011;
        159: y = 16'b1100010100110110;
        160: y = 16'b1100010010001101;
        161: y = 16'b1100001111101110;
        162: y = 16'b1100001101011011;
        163: y = 16'b1100001011010011;
        164: y = 16'b1100001001010110;
        165: y = 16'b1100000111100101;
        166: y = 16'b1100000110000000;
        167: y = 16'b1100000100100111;
        168: y = 16'b1100000011011001;
        169: y = 16'b1100000010010111;
        170: y = 16'b1100000001100001;
        171: y = 16'b1100000000110111;
        172: y = 16'b1100000000011001;
        173: y = 16'b1100000000000111;
        174: y = 16'b1100000000000001;
        175: y = 16'b1100000000000111;
        176: y = 16'b1100000000011001;
        177: y = 16'b1100000000110111;
        178: y = 16'b1100000001100001;
        179: y = 16'b1100000010010111;
        180: y = 16'b1100000011011001;
        181: y = 16'b1100000100100111;
        182: y = 16'b1100000110000000;
        183: y = 16'b1100000111100101;
        184: y = 16'b1100001001010110;
        185: y = 16'b1100001011010011;
        186: y = 16'b1100001101011011;
        187: y = 16'b1100001111101110;
        188: y = 16'b1100010010001101;
        189: y = 16'b1100010100110110;
        190: y = 16'b1100010111101011;
        191: y = 16'b1100011010101011;
        192: y = 16'b1100011101110101;
        193: y = 16'b1100100001001011;
        194: y = 16'b1100100100101010;
        195: y = 16'b1100101000010100;
        196: y = 16'b1100101100001000;
        197: y = 16'b1100110000000110;
        198: y = 16'b1100110100001110;
        199: y = 16'b1100111000011111;
        200: y = 16'b1100111100111001;
        201: y = 16'b1101000001011101;
        202: y = 16'b1101000110001010;
        203: y = 16'b1101001010111111;
        204: y = 16'b1101001111111101;
        205: y = 16'b1101010101000100;
        206: y = 16'b1101011010010010;
        207: y = 16'b1101011111101000;
        208: y = 16'b1101100101000101;
        209: y = 16'b1101101010101010;
        210: y = 16'b1101110000010110;
        211: y = 16'b1101110110001001;
        212: y = 16'b1101111100000010;
        213: y = 16'b1110000010000001;
        214: y = 16'b1110001000000110;
        215: y = 16'b1110001110010001;
        216: y = 16'b1110010100100001;
        217: y = 16'b1110011010110110;
        218: y = 16'b1110100001010000;
        219: y = 16'b1110100111101110;
        220: y = 16'b1110101110010001;
        221: y = 16'b1110110100110111;
        222: y = 16'b1110111011100001;
        223: y = 16'b1111000010001110;
        224: y = 16'b1111001000111110;
        225: y = 16'b1111001111110001;
        226: y = 16'b1111010110100110;
        227: y = 16'b1111011101011100;
        228: y = 16'b1111100100010101;
        229: y = 16'b1111101011001110;
        230: y = 16'b1111110010001001;
        231: y = 16'b1111111001000100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=293.66Hz, Fs=64453Hz, 16-bit

module lut_D
(
    input        [ 7:0] x,
    output       [ 7:0] x_max,
    output logic [15:0] y
);

    assign x_max = 218;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000000111010110;
        2: y = 16'b0000001110101100;
        3: y = 16'b0000010110000000;
        4: y = 16'b0000011101010100;
        5: y = 16'b0000100100100110;
        6: y = 16'b0000101011110110;
        7: y = 16'b0000110011000100;
        8: y = 16'b0000111010001111;
        9: y = 16'b0001000001010111;
        10: y = 16'b0001001000011100;
        11: y = 16'b0001001111011101;
        12: y = 16'b0001010110011010;
        13: y = 16'b0001011101010010;
        14: y = 16'b0001100100000101;
        15: y = 16'b0001101010110011;
        16: y = 16'b0001110001011011;
        17: y = 16'b0001110111111110;
        18: y = 16'b0001111110011010;
        19: y = 16'b0010000100101111;
        20: y = 16'b0010001010111101;
        21: y = 16'b0010010001000100;
        22: y = 16'b0010010111000100;
        23: y = 16'b0010011100111011;
        24: y = 16'b0010100010101010;
        25: y = 16'b0010101000010001;
        26: y = 16'b0010101101101111;
        27: y = 16'b0010110011000011;
        28: y = 16'b0010111000001110;
        29: y = 16'b0010111101010000;
        30: y = 16'b0011000010000111;
        31: y = 16'b0011000110110101;
        32: y = 16'b0011001011010111;
        33: y = 16'b0011001111101111;
        34: y = 16'b0011010011111101;
        35: y = 16'b0011010111111111;
        36: y = 16'b0011011011110101;
        37: y = 16'b0011011111100000;
        38: y = 16'b0011100010111111;
        39: y = 16'b0011100110010011;
        40: y = 16'b0011101001011010;
        41: y = 16'b0011101100010101;
        42: y = 16'b0011101111000011;
        43: y = 16'b0011110001100101;
        44: y = 16'b0011110011111010;
        45: y = 16'b0011110110000010;
        46: y = 16'b0011110111111101;
        47: y = 16'b0011111001101100;
        48: y = 16'b0011111011001101;
        49: y = 16'b0011111100100001;
        50: y = 16'b0011111101100111;
        51: y = 16'b0011111110100000;
        52: y = 16'b0011111111001100;
        53: y = 16'b0011111111101010;
        54: y = 16'b0011111111111011;
        55: y = 16'b0011111111111111;
        56: y = 16'b0011111111110100;
        57: y = 16'b0011111111011101;
        58: y = 16'b0011111110111000;
        59: y = 16'b0011111110000101;
        60: y = 16'b0011111101000110;
        61: y = 16'b0011111011111000;
        62: y = 16'b0011111010011110;
        63: y = 16'b0011111000110110;
        64: y = 16'b0011110111000001;
        65: y = 16'b0011110101000000;
        66: y = 16'b0011110010110001;
        67: y = 16'b0011110000010110;
        68: y = 16'b0011101101101101;
        69: y = 16'b0011101010111001;
        70: y = 16'b0011100111111000;
        71: y = 16'b0011100100101011;
        72: y = 16'b0011100001010001;
        73: y = 16'b0011011101101100;
        74: y = 16'b0011011001111011;
        75: y = 16'b0011010101111111;
        76: y = 16'b0011010001110111;
        77: y = 16'b0011001101100101;
        78: y = 16'b0011001001000111;
        79: y = 16'b0011000100011111;
        80: y = 16'b0010111111101101;
        81: y = 16'b0010111010110000;
        82: y = 16'b0010110101101010;
        83: y = 16'b0010110000011010;
        84: y = 16'b0010101011000001;
        85: y = 16'b0010100101011111;
        86: y = 16'b0010011111110100;
        87: y = 16'b0010011010000000;
        88: y = 16'b0010010100000101;
        89: y = 16'b0010001110000010;
        90: y = 16'b0010000111110111;
        91: y = 16'b0010000001100101;
        92: y = 16'b0001111011001100;
        93: y = 16'b0001110100101101;
        94: y = 16'b0001101110001000;
        95: y = 16'b0001100111011101;
        96: y = 16'b0001100000101100;
        97: y = 16'b0001011001110110;
        98: y = 16'b0001010010111100;
        99: y = 16'b0001001011111101;
        100: y = 16'b0001000100111010;
        101: y = 16'b0000111101110100;
        102: y = 16'b0000110110101010;
        103: y = 16'b0000101111011110;
        104: y = 16'b0000101000001110;
        105: y = 16'b0000100000111101;
        106: y = 16'b0000011001101010;
        107: y = 16'b0000010010010110;
        108: y = 16'b0000001011000001;
        109: y = 16'b0000000011101011;
        110: y = 16'b1111111100010101;
        111: y = 16'b1111110100111111;
        112: y = 16'b1111101101101010;
        113: y = 16'b1111100110010110;
        114: y = 16'b1111011111000011;
        115: y = 16'b1111010111110010;
        116: y = 16'b1111010000100010;
        117: y = 16'b1111001001010110;
        118: y = 16'b1111000010001100;
        119: y = 16'b1110111011000110;
        120: y = 16'b1110110100000011;
        121: y = 16'b1110101101000100;
        122: y = 16'b1110100110001010;
        123: y = 16'b1110011111010100;
        124: y = 16'b1110011000100011;
        125: y = 16'b1110010001111000;
        126: y = 16'b1110001011010011;
        127: y = 16'b1110000100110100;
        128: y = 16'b1101111110011011;
        129: y = 16'b1101111000001001;
        130: y = 16'b1101110001111110;
        131: y = 16'b1101101011111011;
        132: y = 16'b1101100110000000;
        133: y = 16'b1101100000001100;
        134: y = 16'b1101011010100001;
        135: y = 16'b1101010100111111;
        136: y = 16'b1101001111100110;
        137: y = 16'b1101001010010110;
        138: y = 16'b1101000101010000;
        139: y = 16'b1101000000010011;
        140: y = 16'b1100111011100001;
        141: y = 16'b1100110110111001;
        142: y = 16'b1100110010011011;
        143: y = 16'b1100101110001001;
        144: y = 16'b1100101010000001;
        145: y = 16'b1100100110000101;
        146: y = 16'b1100100010010100;
        147: y = 16'b1100011110101111;
        148: y = 16'b1100011011010101;
        149: y = 16'b1100011000001000;
        150: y = 16'b1100010101000111;
        151: y = 16'b1100010010010011;
        152: y = 16'b1100001111101010;
        153: y = 16'b1100001101001111;
        154: y = 16'b1100001011000000;
        155: y = 16'b1100001000111111;
        156: y = 16'b1100000111001010;
        157: y = 16'b1100000101100010;
        158: y = 16'b1100000100001000;
        159: y = 16'b1100000010111010;
        160: y = 16'b1100000001111011;
        161: y = 16'b1100000001001000;
        162: y = 16'b1100000000100011;
        163: y = 16'b1100000000001100;
        164: y = 16'b1100000000000001;
        165: y = 16'b1100000000000101;
        166: y = 16'b1100000000010110;
        167: y = 16'b1100000000110100;
        168: y = 16'b1100000001100000;
        169: y = 16'b1100000010011001;
        170: y = 16'b1100000011011111;
        171: y = 16'b1100000100110011;
        172: y = 16'b1100000110010100;
        173: y = 16'b1100001000000011;
        174: y = 16'b1100001001111110;
        175: y = 16'b1100001100000110;
        176: y = 16'b1100001110011011;
        177: y = 16'b1100010000111101;
        178: y = 16'b1100010011101011;
        179: y = 16'b1100010110100110;
        180: y = 16'b1100011001101101;
        181: y = 16'b1100011101000001;
        182: y = 16'b1100100000100000;
        183: y = 16'b1100100100001011;
        184: y = 16'b1100101000000001;
        185: y = 16'b1100101100000011;
        186: y = 16'b1100110000010001;
        187: y = 16'b1100110100101001;
        188: y = 16'b1100111001001011;
        189: y = 16'b1100111101111001;
        190: y = 16'b1101000010110000;
        191: y = 16'b1101000111110010;
        192: y = 16'b1101001100111101;
        193: y = 16'b1101010010010001;
        194: y = 16'b1101010111101111;
        195: y = 16'b1101011101010110;
        196: y = 16'b1101100011000101;
        197: y = 16'b1101101000111100;
        198: y = 16'b1101101110111100;
        199: y = 16'b1101110101000011;
        200: y = 16'b1101111011010001;
        201: y = 16'b1110000001100110;
        202: y = 16'b1110001000000010;
        203: y = 16'b1110001110100101;
        204: y = 16'b1110010101001101;
        205: y = 16'b1110011011111011;
        206: y = 16'b1110100010101110;
        207: y = 16'b1110101001100110;
        208: y = 16'b1110110000100011;
        209: y = 16'b1110110111100100;
        210: y = 16'b1110111110101001;
        211: y = 16'b1111000101110001;
        212: y = 16'b1111001100111100;
        213: y = 16'b1111010100001010;
        214: y = 16'b1111011011011010;
        215: y = 16'b1111100010101100;
        216: y = 16'b1111101010000000;
        217: y = 16'b1111110001010100;
        218: y = 16'b1111111000101010;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=311.13Hz, Fs=64453Hz, 16-bit

module lut_Ds
(
    input        [ 7:0] x,
    output       [ 7:0] x_max,
    output logic [15:0] y
);

    assign x_max = 206;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000000111110001;
        2: y = 16'b0000001111100010;
        3: y = 16'b0000010111010010;
        4: y = 16'b0000011111000000;
        5: y = 16'b0000100110101101;
        6: y = 16'b0000101110010111;
        7: y = 16'b0000110101111111;
        8: y = 16'b0000111101100011;
        9: y = 16'b0001000101000100;
        10: y = 16'b0001001100100001;
        11: y = 16'b0001010011111001;
        12: y = 16'b0001011011001100;
        13: y = 16'b0001100010011010;
        14: y = 16'b0001101001100010;
        15: y = 16'b0001110000100100;
        16: y = 16'b0001110111011111;
        17: y = 16'b0001111110010100;
        18: y = 16'b0010000101000000;
        19: y = 16'b0010001011100101;
        20: y = 16'b0010010010000010;
        21: y = 16'b0010011000010110;
        22: y = 16'b0010011110100001;
        23: y = 16'b0010100100100011;
        24: y = 16'b0010101010011011;
        25: y = 16'b0010110000001001;
        26: y = 16'b0010110101101100;
        27: y = 16'b0010111011000101;
        28: y = 16'b0011000000010011;
        29: y = 16'b0011000101010110;
        30: y = 16'b0011001010001101;
        31: y = 16'b0011001110110111;
        32: y = 16'b0011010011010110;
        33: y = 16'b0011010111101001;
        34: y = 16'b0011011011101110;
        35: y = 16'b0011011111100111;
        36: y = 16'b0011100011010010;
        37: y = 16'b0011100110110000;
        38: y = 16'b0011101010000001;
        39: y = 16'b0011101101000011;
        40: y = 16'b0011101111111000;
        41: y = 16'b0011110010011111;
        42: y = 16'b0011110100110111;
        43: y = 16'b0011110111000001;
        44: y = 16'b0011111000111100;
        45: y = 16'b0011111010101000;
        46: y = 16'b0011111100000110;
        47: y = 16'b0011111101010101;
        48: y = 16'b0011111110010101;
        49: y = 16'b0011111111000110;
        50: y = 16'b0011111111101000;
        51: y = 16'b0011111111111011;
        52: y = 16'b0011111111111111;
        53: y = 16'b0011111111110011;
        54: y = 16'b0011111111011001;
        55: y = 16'b0011111110101111;
        56: y = 16'b0011111101110111;
        57: y = 16'b0011111100101111;
        58: y = 16'b0011111011011001;
        59: y = 16'b0011111001110100;
        60: y = 16'b0011111000000000;
        61: y = 16'b0011110101111101;
        62: y = 16'b0011110011101100;
        63: y = 16'b0011110001001101;
        64: y = 16'b0011101110011111;
        65: y = 16'b0011101011100100;
        66: y = 16'b0011101000011010;
        67: y = 16'b0011100101000011;
        68: y = 16'b0011100001011110;
        69: y = 16'b0011011101101100;
        70: y = 16'b0011011001101101;
        71: y = 16'b0011010101100001;
        72: y = 16'b0011010001001000;
        73: y = 16'b0011001100100100;
        74: y = 16'b0011000111110011;
        75: y = 16'b0011000010110110;
        76: y = 16'b0010111101101110;
        77: y = 16'b0010111000011010;
        78: y = 16'b0010110010111100;
        79: y = 16'b0010101101010011;
        80: y = 16'b0010100111100000;
        81: y = 16'b0010100001100011;
        82: y = 16'b0010011011011101;
        83: y = 16'b0010010101001101;
        84: y = 16'b0010001110110101;
        85: y = 16'b0010001000010100;
        86: y = 16'b0010000001101011;
        87: y = 16'b0001111010111010;
        88: y = 16'b0001110100000011;
        89: y = 16'b0001101101000100;
        90: y = 16'b0001100101111111;
        91: y = 16'b0001011110110100;
        92: y = 16'b0001010111100011;
        93: y = 16'b0001010000001110;
        94: y = 16'b0001001000110011;
        95: y = 16'b0001000001010100;
        96: y = 16'b0000111001110001;
        97: y = 16'b0000110010001011;
        98: y = 16'b0000101010100010;
        99: y = 16'b0000100010110111;
        100: y = 16'b0000011011001001;
        101: y = 16'b0000010011011010;
        102: y = 16'b0000001011101010;
        103: y = 16'b0000000011111001;
        104: y = 16'b1111111100000111;
        105: y = 16'b1111110100010110;
        106: y = 16'b1111101100100110;
        107: y = 16'b1111100100110111;
        108: y = 16'b1111011101001001;
        109: y = 16'b1111010101011110;
        110: y = 16'b1111001101110101;
        111: y = 16'b1111000110001111;
        112: y = 16'b1110111110101100;
        113: y = 16'b1110110111001101;
        114: y = 16'b1110101111110010;
        115: y = 16'b1110101000011101;
        116: y = 16'b1110100001001100;
        117: y = 16'b1110011010000001;
        118: y = 16'b1110010010111100;
        119: y = 16'b1110001011111101;
        120: y = 16'b1110000101000110;
        121: y = 16'b1101111110010101;
        122: y = 16'b1101110111101100;
        123: y = 16'b1101110001001011;
        124: y = 16'b1101101010110011;
        125: y = 16'b1101100100100011;
        126: y = 16'b1101011110011101;
        127: y = 16'b1101011000100000;
        128: y = 16'b1101010010101101;
        129: y = 16'b1101001101000100;
        130: y = 16'b1101000111100110;
        131: y = 16'b1101000010010010;
        132: y = 16'b1100111101001010;
        133: y = 16'b1100111000001101;
        134: y = 16'b1100110011011100;
        135: y = 16'b1100101110111000;
        136: y = 16'b1100101010011111;
        137: y = 16'b1100100110010011;
        138: y = 16'b1100100010010100;
        139: y = 16'b1100011110100010;
        140: y = 16'b1100011010111101;
        141: y = 16'b1100010111100110;
        142: y = 16'b1100010100011100;
        143: y = 16'b1100010001100001;
        144: y = 16'b1100001110110011;
        145: y = 16'b1100001100010100;
        146: y = 16'b1100001010000011;
        147: y = 16'b1100001000000000;
        148: y = 16'b1100000110001100;
        149: y = 16'b1100000100100111;
        150: y = 16'b1100000011010001;
        151: y = 16'b1100000010001001;
        152: y = 16'b1100000001010001;
        153: y = 16'b1100000000100111;
        154: y = 16'b1100000000001101;
        155: y = 16'b1100000000000001;
        156: y = 16'b1100000000000101;
        157: y = 16'b1100000000011000;
        158: y = 16'b1100000000111010;
        159: y = 16'b1100000001101011;
        160: y = 16'b1100000010101011;
        161: y = 16'b1100000011111010;
        162: y = 16'b1100000101011000;
        163: y = 16'b1100000111000100;
        164: y = 16'b1100001000111111;
        165: y = 16'b1100001011001001;
        166: y = 16'b1100001101100001;
        167: y = 16'b1100010000001000;
        168: y = 16'b1100010010111101;
        169: y = 16'b1100010101111111;
        170: y = 16'b1100011001010000;
        171: y = 16'b1100011100101110;
        172: y = 16'b1100100000011001;
        173: y = 16'b1100100100010010;
        174: y = 16'b1100101000010111;
        175: y = 16'b1100101100101010;
        176: y = 16'b1100110001001001;
        177: y = 16'b1100110101110011;
        178: y = 16'b1100111010101010;
        179: y = 16'b1100111111101101;
        180: y = 16'b1101000100111011;
        181: y = 16'b1101001010010100;
        182: y = 16'b1101001111110111;
        183: y = 16'b1101010101100101;
        184: y = 16'b1101011011011101;
        185: y = 16'b1101100001011111;
        186: y = 16'b1101100111101010;
        187: y = 16'b1101101101111110;
        188: y = 16'b1101110100011011;
        189: y = 16'b1101111011000000;
        190: y = 16'b1110000001101100;
        191: y = 16'b1110001000100001;
        192: y = 16'b1110001111011100;
        193: y = 16'b1110010110011110;
        194: y = 16'b1110011101100110;
        195: y = 16'b1110100100110100;
        196: y = 16'b1110101100000111;
        197: y = 16'b1110110011011111;
        198: y = 16'b1110111010111100;
        199: y = 16'b1111000010011101;
        200: y = 16'b1111001010000001;
        201: y = 16'b1111010001101001;
        202: y = 16'b1111011001010011;
        203: y = 16'b1111100001000000;
        204: y = 16'b1111101000101110;
        205: y = 16'b1111110000011110;
        206: y = 16'b1111111000001111;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=329.63Hz, Fs=64453Hz, 16-bit

module lut_E
(
    input        [ 7:0] x,
    output       [ 7:0] x_max,
    output logic [15:0] y
);

    assign x_max = 194;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001000010000;
        2: y = 16'b0000010000011111;
        3: y = 16'b0000011000101101;
        4: y = 16'b0000100000111010;
        5: y = 16'b0000101001000100;
        6: y = 16'b0000110001001100;
        7: y = 16'b0000111001010000;
        8: y = 16'b0001000001010000;
        9: y = 16'b0001001001001101;
        10: y = 16'b0001010001000100;
        11: y = 16'b0001011000110110;
        12: y = 16'b0001100000100010;
        13: y = 16'b0001101000001000;
        14: y = 16'b0001101111100110;
        15: y = 16'b0001110110111110;
        16: y = 16'b0001111110001101;
        17: y = 16'b0010000101010100;
        18: y = 16'b0010001100010010;
        19: y = 16'b0010010011000111;
        20: y = 16'b0010011001110010;
        21: y = 16'b0010100000010011;
        22: y = 16'b0010100110101001;
        23: y = 16'b0010101100110100;
        24: y = 16'b0010110010110100;
        25: y = 16'b0010111000100111;
        26: y = 16'b0010111110001111;
        27: y = 16'b0011000011101010;
        28: y = 16'b0011001000111000;
        29: y = 16'b0011001101111000;
        30: y = 16'b0011010010101011;
        31: y = 16'b0011010111010000;
        32: y = 16'b0011011011100110;
        33: y = 16'b0011011111101110;
        34: y = 16'b0011100011100111;
        35: y = 16'b0011100111010001;
        36: y = 16'b0011101010101100;
        37: y = 16'b0011101101110111;
        38: y = 16'b0011110000110010;
        39: y = 16'b0011110011011101;
        40: y = 16'b0011110101111000;
        41: y = 16'b0011111000000011;
        42: y = 16'b0011111001111101;
        43: y = 16'b0011111011100111;
        44: y = 16'b0011111100111111;
        45: y = 16'b0011111110001000;
        46: y = 16'b0011111110111111;
        47: y = 16'b0011111111100101;
        48: y = 16'b0011111111111010;
        49: y = 16'b0011111111111110;
        50: y = 16'b0011111111110010;
        51: y = 16'b0011111111010100;
        52: y = 16'b0011111110100101;
        53: y = 16'b0011111101100110;
        54: y = 16'b0011111100010101;
        55: y = 16'b0011111010110100;
        56: y = 16'b0011111001000010;
        57: y = 16'b0011110111000000;
        58: y = 16'b0011110100101101;
        59: y = 16'b0011110010001010;
        60: y = 16'b0011101111010110;
        61: y = 16'b0011101100010011;
        62: y = 16'b0011101001000000;
        63: y = 16'b0011100101011110;
        64: y = 16'b0011100001101101;
        65: y = 16'b0011011101101100;
        66: y = 16'b0011011001011101;
        67: y = 16'b0011010100111111;
        68: y = 16'b0011010000010011;
        69: y = 16'b0011001011011010;
        70: y = 16'b0011000110010010;
        71: y = 16'b0011000000111110;
        72: y = 16'b0010111011011101;
        73: y = 16'b0010110101101111;
        74: y = 16'b0010101111110101;
        75: y = 16'b0010101001110000;
        76: y = 16'b0010100011011111;
        77: y = 16'b0010011101000100;
        78: y = 16'b0010010110011110;
        79: y = 16'b0010001111101110;
        80: y = 16'b0010001000110100;
        81: y = 16'b0010000001110010;
        82: y = 16'b0001111010100110;
        83: y = 16'b0001110011010011;
        84: y = 16'b0001101011111000;
        85: y = 16'b0001100100010110;
        86: y = 16'b0001011100101101;
        87: y = 16'b0001010100111110;
        88: y = 16'b0001001101001001;
        89: y = 16'b0001000101001111;
        90: y = 16'b0000111101010001;
        91: y = 16'b0000110101001110;
        92: y = 16'b0000101101001000;
        93: y = 16'b0000100100111111;
        94: y = 16'b0000011100110100;
        95: y = 16'b0000010100100110;
        96: y = 16'b0000001100011000;
        97: y = 16'b0000000100001000;
        98: y = 16'b1111111011111000;
        99: y = 16'b1111110011101000;
        100: y = 16'b1111101011011010;
        101: y = 16'b1111100011001100;
        102: y = 16'b1111011011000001;
        103: y = 16'b1111010010111000;
        104: y = 16'b1111001010110010;
        105: y = 16'b1111000010101111;
        106: y = 16'b1110111010110001;
        107: y = 16'b1110110010110111;
        108: y = 16'b1110101011000010;
        109: y = 16'b1110100011010011;
        110: y = 16'b1110011011101010;
        111: y = 16'b1110010100001000;
        112: y = 16'b1110001100101101;
        113: y = 16'b1110000101011010;
        114: y = 16'b1101111110001110;
        115: y = 16'b1101110111001100;
        116: y = 16'b1101110000010010;
        117: y = 16'b1101101001100010;
        118: y = 16'b1101100010111100;
        119: y = 16'b1101011100100001;
        120: y = 16'b1101010110010000;
        121: y = 16'b1101010000001011;
        122: y = 16'b1101001010010001;
        123: y = 16'b1101000100100011;
        124: y = 16'b1100111111000010;
        125: y = 16'b1100111001101110;
        126: y = 16'b1100110100100110;
        127: y = 16'b1100101111101101;
        128: y = 16'b1100101011000001;
        129: y = 16'b1100100110100011;
        130: y = 16'b1100100010010100;
        131: y = 16'b1100011110010011;
        132: y = 16'b1100011010100010;
        133: y = 16'b1100010111000000;
        134: y = 16'b1100010011101101;
        135: y = 16'b1100010000101010;
        136: y = 16'b1100001101110110;
        137: y = 16'b1100001011010011;
        138: y = 16'b1100001001000000;
        139: y = 16'b1100000110111110;
        140: y = 16'b1100000101001100;
        141: y = 16'b1100000011101011;
        142: y = 16'b1100000010011010;
        143: y = 16'b1100000001011011;
        144: y = 16'b1100000000101100;
        145: y = 16'b1100000000001110;
        146: y = 16'b1100000000000010;
        147: y = 16'b1100000000000110;
        148: y = 16'b1100000000011011;
        149: y = 16'b1100000001000001;
        150: y = 16'b1100000001111000;
        151: y = 16'b1100000011000001;
        152: y = 16'b1100000100011001;
        153: y = 16'b1100000110000011;
        154: y = 16'b1100000111111101;
        155: y = 16'b1100001010001000;
        156: y = 16'b1100001100100011;
        157: y = 16'b1100001111001110;
        158: y = 16'b1100010010001001;
        159: y = 16'b1100010101010100;
        160: y = 16'b1100011000101111;
        161: y = 16'b1100011100011001;
        162: y = 16'b1100100000010010;
        163: y = 16'b1100100100011010;
        164: y = 16'b1100101000110000;
        165: y = 16'b1100101101010101;
        166: y = 16'b1100110010001000;
        167: y = 16'b1100110111001000;
        168: y = 16'b1100111100010110;
        169: y = 16'b1101000001110001;
        170: y = 16'b1101000111011001;
        171: y = 16'b1101001101001100;
        172: y = 16'b1101010011001100;
        173: y = 16'b1101011001010111;
        174: y = 16'b1101011111101101;
        175: y = 16'b1101100110001110;
        176: y = 16'b1101101100111001;
        177: y = 16'b1101110011101110;
        178: y = 16'b1101111010101100;
        179: y = 16'b1110000001110011;
        180: y = 16'b1110001001000010;
        181: y = 16'b1110010000011010;
        182: y = 16'b1110010111111000;
        183: y = 16'b1110011111011110;
        184: y = 16'b1110100111001010;
        185: y = 16'b1110101110111100;
        186: y = 16'b1110110110110011;
        187: y = 16'b1110111110110000;
        188: y = 16'b1111000110110000;
        189: y = 16'b1111001110110100;
        190: y = 16'b1111010110111100;
        191: y = 16'b1111011111000110;
        192: y = 16'b1111100111010011;
        193: y = 16'b1111101111100001;
        194: y = 16'b1111110111110000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=349.23Hz, Fs=64453Hz, 16-bit

module lut_F
(
    input        [ 7:0] x,
    output       [ 7:0] x_max,
    output logic [15:0] y
);

    assign x_max = 183;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001000101111;
        2: y = 16'b0000010001011110;
        3: y = 16'b0000011010001011;
        4: y = 16'b0000100010110111;
        5: y = 16'b0000101011100000;
        6: y = 16'b0000110100000101;
        7: y = 16'b0000111100100111;
        8: y = 16'b0001000101000100;
        9: y = 16'b0001001101011100;
        10: y = 16'b0001010101101110;
        11: y = 16'b0001011101111010;
        12: y = 16'b0001100101111111;
        13: y = 16'b0001101101111100;
        14: y = 16'b0001110101110001;
        15: y = 16'b0001111101011101;
        16: y = 16'b0010000101000000;
        17: y = 16'b0010001100011001;
        18: y = 16'b0010010011101000;
        19: y = 16'b0010011010101011;
        20: y = 16'b0010100001100011;
        21: y = 16'b0010101000001111;
        22: y = 16'b0010101110101110;
        23: y = 16'b0010110101000001;
        24: y = 16'b0010111011000101;
        25: y = 16'b0011000000111100;
        26: y = 16'b0011000110100100;
        27: y = 16'b0011001011111110;
        28: y = 16'b0011010001001000;
        29: y = 16'b0011010110000011;
        30: y = 16'b0011011010101110;
        31: y = 16'b0011011111001000;
        32: y = 16'b0011100011010010;
        33: y = 16'b0011100111001011;
        34: y = 16'b0011101010110011;
        35: y = 16'b0011101110001001;
        36: y = 16'b0011110001001101;
        37: y = 16'b0011110011111111;
        38: y = 16'b0011110110011111;
        39: y = 16'b0011111000101101;
        40: y = 16'b0011111010101000;
        41: y = 16'b0011111100010001;
        42: y = 16'b0011111101100110;
        43: y = 16'b0011111110101001;
        44: y = 16'b0011111111011001;
        45: y = 16'b0011111111110101;
        46: y = 16'b0011111111111111;
        47: y = 16'b0011111111110101;
        48: y = 16'b0011111111011001;
        49: y = 16'b0011111110101001;
        50: y = 16'b0011111101100110;
        51: y = 16'b0011111100010001;
        52: y = 16'b0011111010101000;
        53: y = 16'b0011111000101101;
        54: y = 16'b0011110110011111;
        55: y = 16'b0011110011111111;
        56: y = 16'b0011110001001101;
        57: y = 16'b0011101110001001;
        58: y = 16'b0011101010110011;
        59: y = 16'b0011100111001011;
        60: y = 16'b0011100011010010;
        61: y = 16'b0011011111001000;
        62: y = 16'b0011011010101110;
        63: y = 16'b0011010110000011;
        64: y = 16'b0011010001001000;
        65: y = 16'b0011001011111110;
        66: y = 16'b0011000110100100;
        67: y = 16'b0011000000111100;
        68: y = 16'b0010111011000101;
        69: y = 16'b0010110101000001;
        70: y = 16'b0010101110101110;
        71: y = 16'b0010101000001111;
        72: y = 16'b0010100001100011;
        73: y = 16'b0010011010101011;
        74: y = 16'b0010010011101000;
        75: y = 16'b0010001100011001;
        76: y = 16'b0010000101000000;
        77: y = 16'b0001111101011101;
        78: y = 16'b0001110101110001;
        79: y = 16'b0001101101111100;
        80: y = 16'b0001100101111111;
        81: y = 16'b0001011101111010;
        82: y = 16'b0001010101101110;
        83: y = 16'b0001001101011100;
        84: y = 16'b0001000101000100;
        85: y = 16'b0000111100100111;
        86: y = 16'b0000110100000101;
        87: y = 16'b0000101011100000;
        88: y = 16'b0000100010110111;
        89: y = 16'b0000011010001011;
        90: y = 16'b0000010001011110;
        91: y = 16'b0000001000101111;
        92: y = 16'b0000000000000000;
        93: y = 16'b1111110111010001;
        94: y = 16'b1111101110100010;
        95: y = 16'b1111100101110101;
        96: y = 16'b1111011101001001;
        97: y = 16'b1111010100100000;
        98: y = 16'b1111001011111011;
        99: y = 16'b1111000011011001;
        100: y = 16'b1110111010111100;
        101: y = 16'b1110110010100100;
        102: y = 16'b1110101010010010;
        103: y = 16'b1110100010000110;
        104: y = 16'b1110011010000001;
        105: y = 16'b1110010010000100;
        106: y = 16'b1110001010001111;
        107: y = 16'b1110000010100011;
        108: y = 16'b1101111011000000;
        109: y = 16'b1101110011100111;
        110: y = 16'b1101101100011000;
        111: y = 16'b1101100101010101;
        112: y = 16'b1101011110011101;
        113: y = 16'b1101010111110001;
        114: y = 16'b1101010001010010;
        115: y = 16'b1101001010111111;
        116: y = 16'b1101000100111011;
        117: y = 16'b1100111111000100;
        118: y = 16'b1100111001011100;
        119: y = 16'b1100110100000010;
        120: y = 16'b1100101110111000;
        121: y = 16'b1100101001111101;
        122: y = 16'b1100100101010010;
        123: y = 16'b1100100000111000;
        124: y = 16'b1100011100101110;
        125: y = 16'b1100011000110101;
        126: y = 16'b1100010101001101;
        127: y = 16'b1100010001110111;
        128: y = 16'b1100001110110011;
        129: y = 16'b1100001100000001;
        130: y = 16'b1100001001100001;
        131: y = 16'b1100000111010011;
        132: y = 16'b1100000101011000;
        133: y = 16'b1100000011101111;
        134: y = 16'b1100000010011010;
        135: y = 16'b1100000001010111;
        136: y = 16'b1100000000100111;
        137: y = 16'b1100000000001011;
        138: y = 16'b1100000000000001;
        139: y = 16'b1100000000001011;
        140: y = 16'b1100000000100111;
        141: y = 16'b1100000001010111;
        142: y = 16'b1100000010011010;
        143: y = 16'b1100000011101111;
        144: y = 16'b1100000101011000;
        145: y = 16'b1100000111010011;
        146: y = 16'b1100001001100001;
        147: y = 16'b1100001100000001;
        148: y = 16'b1100001110110011;
        149: y = 16'b1100010001110111;
        150: y = 16'b1100010101001101;
        151: y = 16'b1100011000110101;
        152: y = 16'b1100011100101110;
        153: y = 16'b1100100000111000;
        154: y = 16'b1100100101010010;
        155: y = 16'b1100101001111101;
        156: y = 16'b1100101110111000;
        157: y = 16'b1100110100000010;
        158: y = 16'b1100111001011100;
        159: y = 16'b1100111111000100;
        160: y = 16'b1101000100111011;
        161: y = 16'b1101001010111111;
        162: y = 16'b1101010001010010;
        163: y = 16'b1101010111110001;
        164: y = 16'b1101011110011101;
        165: y = 16'b1101100101010101;
        166: y = 16'b1101101100011000;
        167: y = 16'b1101110011100111;
        168: y = 16'b1101111011000000;
        169: y = 16'b1110000010100011;
        170: y = 16'b1110001010001111;
        171: y = 16'b1110010010000100;
        172: y = 16'b1110011010000001;
        173: y = 16'b1110100010000110;
        174: y = 16'b1110101010010010;
        175: y = 16'b1110110010100100;
        176: y = 16'b1110111010111100;
        177: y = 16'b1111000011011001;
        178: y = 16'b1111001011111011;
        179: y = 16'b1111010100100000;
        180: y = 16'b1111011101001001;
        181: y = 16'b1111100101110101;
        182: y = 16'b1111101110100010;
        183: y = 16'b1111110111010001;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=369.99Hz, Fs=64453Hz, 16-bit

module lut_Fs
(
    input        [ 7:0] x,
    output       [ 7:0] x_max,
    output logic [15:0] y
);

    assign x_max = 173;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001001001111;
        2: y = 16'b0000010010011110;
        3: y = 16'b0000011011101011;
        4: y = 16'b0000100100110110;
        5: y = 16'b0000101101111110;
        6: y = 16'b0000110111000010;
        7: y = 16'b0001000000000001;
        8: y = 16'b0001001000111011;
        9: y = 16'b0001010001101111;
        10: y = 16'b0001011010011100;
        11: y = 16'b0001100011000010;
        12: y = 16'b0001101011011111;
        13: y = 16'b0001110011110011;
        14: y = 16'b0001111011111110;
        15: y = 16'b0010000011111110;
        16: y = 16'b0010001011110100;
        17: y = 16'b0010010011011101;
        18: y = 16'b0010011010111011;
        19: y = 16'b0010100010001011;
        20: y = 16'b0010101001001110;
        21: y = 16'b0010110000000011;
        22: y = 16'b0010110110101001;
        23: y = 16'b0010111100111111;
        24: y = 16'b0011000011000111;
        25: y = 16'b0011001000111101;
        26: y = 16'b0011001110100011;
        27: y = 16'b0011010011111000;
        28: y = 16'b0011011000111011;
        29: y = 16'b0011011101101100;
        30: y = 16'b0011100010001011;
        31: y = 16'b0011100110010110;
        32: y = 16'b0011101010001111;
        33: y = 16'b0011101101110011;
        34: y = 16'b0011110001000100;
        35: y = 16'b0011110100000001;
        36: y = 16'b0011110110101010;
        37: y = 16'b0011111000111110;
        38: y = 16'b0011111010111101;
        39: y = 16'b0011111100100111;
        40: y = 16'b0011111101111100;
        41: y = 16'b0011111110111100;
        42: y = 16'b0011111111100111;
        43: y = 16'b0011111111111100;
        44: y = 16'b0011111111111100;
        45: y = 16'b0011111111100111;
        46: y = 16'b0011111110111100;
        47: y = 16'b0011111101111100;
        48: y = 16'b0011111100100111;
        49: y = 16'b0011111010111101;
        50: y = 16'b0011111000111110;
        51: y = 16'b0011110110101010;
        52: y = 16'b0011110100000001;
        53: y = 16'b0011110001000100;
        54: y = 16'b0011101101110011;
        55: y = 16'b0011101010001111;
        56: y = 16'b0011100110010110;
        57: y = 16'b0011100010001011;
        58: y = 16'b0011011101101100;
        59: y = 16'b0011011000111011;
        60: y = 16'b0011010011111000;
        61: y = 16'b0011001110100011;
        62: y = 16'b0011001000111101;
        63: y = 16'b0011000011000111;
        64: y = 16'b0010111100111111;
        65: y = 16'b0010110110101001;
        66: y = 16'b0010110000000011;
        67: y = 16'b0010101001001110;
        68: y = 16'b0010100010001011;
        69: y = 16'b0010011010111011;
        70: y = 16'b0010010011011101;
        71: y = 16'b0010001011110100;
        72: y = 16'b0010000011111110;
        73: y = 16'b0001111011111110;
        74: y = 16'b0001110011110011;
        75: y = 16'b0001101011011111;
        76: y = 16'b0001100011000010;
        77: y = 16'b0001011010011100;
        78: y = 16'b0001010001101111;
        79: y = 16'b0001001000111011;
        80: y = 16'b0001000000000001;
        81: y = 16'b0000110111000010;
        82: y = 16'b0000101101111110;
        83: y = 16'b0000100100110110;
        84: y = 16'b0000011011101011;
        85: y = 16'b0000010010011110;
        86: y = 16'b0000001001001111;
        87: y = 16'b0000000000000000;
        88: y = 16'b1111110110110001;
        89: y = 16'b1111101101100010;
        90: y = 16'b1111100100010101;
        91: y = 16'b1111011011001010;
        92: y = 16'b1111010010000010;
        93: y = 16'b1111001000111110;
        94: y = 16'b1110111111111111;
        95: y = 16'b1110110111000101;
        96: y = 16'b1110101110010001;
        97: y = 16'b1110100101100100;
        98: y = 16'b1110011100111110;
        99: y = 16'b1110010100100001;
        100: y = 16'b1110001100001101;
        101: y = 16'b1110000100000010;
        102: y = 16'b1101111100000010;
        103: y = 16'b1101110100001100;
        104: y = 16'b1101101100100011;
        105: y = 16'b1101100101000101;
        106: y = 16'b1101011101110101;
        107: y = 16'b1101010110110010;
        108: y = 16'b1101001111111101;
        109: y = 16'b1101001001010111;
        110: y = 16'b1101000011000001;
        111: y = 16'b1100111100111001;
        112: y = 16'b1100110111000011;
        113: y = 16'b1100110001011101;
        114: y = 16'b1100101100001000;
        115: y = 16'b1100100111000101;
        116: y = 16'b1100100010010100;
        117: y = 16'b1100011101110101;
        118: y = 16'b1100011001101010;
        119: y = 16'b1100010101110001;
        120: y = 16'b1100010010001101;
        121: y = 16'b1100001110111100;
        122: y = 16'b1100001011111111;
        123: y = 16'b1100001001010110;
        124: y = 16'b1100000111000010;
        125: y = 16'b1100000101000011;
        126: y = 16'b1100000011011001;
        127: y = 16'b1100000010000100;
        128: y = 16'b1100000001000100;
        129: y = 16'b1100000000011001;
        130: y = 16'b1100000000000100;
        131: y = 16'b1100000000000100;
        132: y = 16'b1100000000011001;
        133: y = 16'b1100000001000100;
        134: y = 16'b1100000010000100;
        135: y = 16'b1100000011011001;
        136: y = 16'b1100000101000011;
        137: y = 16'b1100000111000010;
        138: y = 16'b1100001001010110;
        139: y = 16'b1100001011111111;
        140: y = 16'b1100001110111100;
        141: y = 16'b1100010010001101;
        142: y = 16'b1100010101110001;
        143: y = 16'b1100011001101010;
        144: y = 16'b1100011101110101;
        145: y = 16'b1100100010010100;
        146: y = 16'b1100100111000101;
        147: y = 16'b1100101100001000;
        148: y = 16'b1100110001011101;
        149: y = 16'b1100110111000011;
        150: y = 16'b1100111100111001;
        151: y = 16'b1101000011000001;
        152: y = 16'b1101001001010111;
        153: y = 16'b1101001111111101;
        154: y = 16'b1101010110110010;
        155: y = 16'b1101011101110101;
        156: y = 16'b1101100101000101;
        157: y = 16'b1101101100100011;
        158: y = 16'b1101110100001100;
        159: y = 16'b1101111100000010;
        160: y = 16'b1110000100000010;
        161: y = 16'b1110001100001101;
        162: y = 16'b1110010100100001;
        163: y = 16'b1110011100111110;
        164: y = 16'b1110100101100100;
        165: y = 16'b1110101110010001;
        166: y = 16'b1110110111000101;
        167: y = 16'b1110111111111111;
        168: y = 16'b1111001000111110;
        169: y = 16'b1111010010000010;
        170: y = 16'b1111011011001010;
        171: y = 16'b1111100100010101;
        172: y = 16'b1111101101100010;
        173: y = 16'b1111110110110001;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=392.0Hz, Fs=64453Hz, 16-bit

module lut_G
(
    input        [ 7:0] x,
    output       [ 7:0] x_max,
    output logic [15:0] y
);

    assign x_max = 163;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001001110100;
        2: y = 16'b0000010011100110;
        3: y = 16'b0000011101010111;
        4: y = 16'b0000100111000101;
        5: y = 16'b0000110000101111;
        6: y = 16'b0000111010010101;
        7: y = 16'b0001000011110101;
        8: y = 16'b0001001101001111;
        9: y = 16'b0001010110100010;
        10: y = 16'b0001011111101100;
        11: y = 16'b0001101000101110;
        12: y = 16'b0001110001100101;
        13: y = 16'b0001111010010010;
        14: y = 16'b0010000010110100;
        15: y = 16'b0010001011001001;
        16: y = 16'b0010010011010001;
        17: y = 16'b0010011011001100;
        18: y = 16'b0010100010111000;
        19: y = 16'b0010101010010100;
        20: y = 16'b0010110001100001;
        21: y = 16'b0010111000011100;
        22: y = 16'b0010111111000111;
        23: y = 16'b0011000101011111;
        24: y = 16'b0011001011100101;
        25: y = 16'b0011010001011000;
        26: y = 16'b0011010110110111;
        27: y = 16'b0011011100000010;
        28: y = 16'b0011100000111001;
        29: y = 16'b0011100101011010;
        30: y = 16'b0011101001100110;
        31: y = 16'b0011101101011011;
        32: y = 16'b0011110000111011;
        33: y = 16'b0011110100000011;
        34: y = 16'b0011110110110101;
        35: y = 16'b0011111001010000;
        36: y = 16'b0011111011010011;
        37: y = 16'b0011111100111111;
        38: y = 16'b0011111110010011;
        39: y = 16'b0011111111001111;
        40: y = 16'b0011111111110011;
        41: y = 16'b0011111111111111;
        42: y = 16'b0011111111110011;
        43: y = 16'b0011111111001111;
        44: y = 16'b0011111110010011;
        45: y = 16'b0011111100111111;
        46: y = 16'b0011111011010011;
        47: y = 16'b0011111001010000;
        48: y = 16'b0011110110110101;
        49: y = 16'b0011110100000011;
        50: y = 16'b0011110000111011;
        51: y = 16'b0011101101011011;
        52: y = 16'b0011101001100110;
        53: y = 16'b0011100101011010;
        54: y = 16'b0011100000111001;
        55: y = 16'b0011011100000010;
        56: y = 16'b0011010110110111;
        57: y = 16'b0011010001011000;
        58: y = 16'b0011001011100101;
        59: y = 16'b0011000101011111;
        60: y = 16'b0010111111000111;
        61: y = 16'b0010111000011100;
        62: y = 16'b0010110001100001;
        63: y = 16'b0010101010010100;
        64: y = 16'b0010100010111000;
        65: y = 16'b0010011011001100;
        66: y = 16'b0010010011010001;
        67: y = 16'b0010001011001001;
        68: y = 16'b0010000010110100;
        69: y = 16'b0001111010010010;
        70: y = 16'b0001110001100101;
        71: y = 16'b0001101000101110;
        72: y = 16'b0001011111101100;
        73: y = 16'b0001010110100010;
        74: y = 16'b0001001101001111;
        75: y = 16'b0001000011110101;
        76: y = 16'b0000111010010101;
        77: y = 16'b0000110000101111;
        78: y = 16'b0000100111000101;
        79: y = 16'b0000011101010111;
        80: y = 16'b0000010011100110;
        81: y = 16'b0000001001110100;
        82: y = 16'b0000000000000000;
        83: y = 16'b1111110110001100;
        84: y = 16'b1111101100011010;
        85: y = 16'b1111100010101001;
        86: y = 16'b1111011000111011;
        87: y = 16'b1111001111010001;
        88: y = 16'b1111000101101011;
        89: y = 16'b1110111100001011;
        90: y = 16'b1110110010110001;
        91: y = 16'b1110101001011110;
        92: y = 16'b1110100000010100;
        93: y = 16'b1110010111010010;
        94: y = 16'b1110001110011011;
        95: y = 16'b1110000101101110;
        96: y = 16'b1101111101001100;
        97: y = 16'b1101110100110111;
        98: y = 16'b1101101100101111;
        99: y = 16'b1101100100110100;
        100: y = 16'b1101011101001000;
        101: y = 16'b1101010101101100;
        102: y = 16'b1101001110011111;
        103: y = 16'b1101000111100100;
        104: y = 16'b1101000000111001;
        105: y = 16'b1100111010100001;
        106: y = 16'b1100110100011011;
        107: y = 16'b1100101110101000;
        108: y = 16'b1100101001001001;
        109: y = 16'b1100100011111110;
        110: y = 16'b1100011111000111;
        111: y = 16'b1100011010100110;
        112: y = 16'b1100010110011010;
        113: y = 16'b1100010010100101;
        114: y = 16'b1100001111000101;
        115: y = 16'b1100001011111101;
        116: y = 16'b1100001001001011;
        117: y = 16'b1100000110110000;
        118: y = 16'b1100000100101101;
        119: y = 16'b1100000011000001;
        120: y = 16'b1100000001101101;
        121: y = 16'b1100000000110001;
        122: y = 16'b1100000000001101;
        123: y = 16'b1100000000000001;
        124: y = 16'b1100000000001101;
        125: y = 16'b1100000000110001;
        126: y = 16'b1100000001101101;
        127: y = 16'b1100000011000001;
        128: y = 16'b1100000100101101;
        129: y = 16'b1100000110110000;
        130: y = 16'b1100001001001011;
        131: y = 16'b1100001011111101;
        132: y = 16'b1100001111000101;
        133: y = 16'b1100010010100101;
        134: y = 16'b1100010110011010;
        135: y = 16'b1100011010100110;
        136: y = 16'b1100011111000111;
        137: y = 16'b1100100011111110;
        138: y = 16'b1100101001001001;
        139: y = 16'b1100101110101000;
        140: y = 16'b1100110100011011;
        141: y = 16'b1100111010100001;
        142: y = 16'b1101000000111001;
        143: y = 16'b1101000111100100;
        144: y = 16'b1101001110011111;
        145: y = 16'b1101010101101100;
        146: y = 16'b1101011101001000;
        147: y = 16'b1101100100110100;
        148: y = 16'b1101101100101111;
        149: y = 16'b1101110100110111;
        150: y = 16'b1101111101001100;
        151: y = 16'b1110000101101110;
        152: y = 16'b1110001110011011;
        153: y = 16'b1110010111010010;
        154: y = 16'b1110100000010100;
        155: y = 16'b1110101001011110;
        156: y = 16'b1110110010110001;
        157: y = 16'b1110111100001011;
        158: y = 16'b1111000101101011;
        159: y = 16'b1111001111010001;
        160: y = 16'b1111011000111011;
        161: y = 16'b1111100010101001;
        162: y = 16'b1111101100011010;
        163: y = 16'b1111110110001100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=415.3Hz, Fs=64453Hz, 16-bit

module lut_Gs
(
    input        [ 7:0] x,
    output       [ 7:0] x_max,
    output logic [15:0] y
);

    assign x_max = 154;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001010011000;
        2: y = 16'b0000010100101111;
        3: y = 16'b0000011111000011;
        4: y = 16'b0000101001010101;
        5: y = 16'b0000110011100010;
        6: y = 16'b0000111101101010;
        7: y = 16'b0001000111101011;
        8: y = 16'b0001010001100100;
        9: y = 16'b0001011011010101;
        10: y = 16'b0001100100111101;
        11: y = 16'b0001101110011010;
        12: y = 16'b0001110111101011;
        13: y = 16'b0010000000101111;
        14: y = 16'b0010001001100110;
        15: y = 16'b0010010010001111;
        16: y = 16'b0010011010101000;
        17: y = 16'b0010100010110001;
        18: y = 16'b0010101010101001;
        19: y = 16'b0010110010001111;
        20: y = 16'b0010111001100010;
        21: y = 16'b0011000000100010;
        22: y = 16'b0011000111001101;
        23: y = 16'b0011001101100100;
        24: y = 16'b0011010011100101;
        25: y = 16'b0011011001001111;
        26: y = 16'b0011011110100011;
        27: y = 16'b0011100011011111;
        28: y = 16'b0011101000000100;
        29: y = 16'b0011101100010000;
        30: y = 16'b0011110000000011;
        31: y = 16'b0011110011011101;
        32: y = 16'b0011110110011110;
        33: y = 16'b0011111001000100;
        34: y = 16'b0011111011010000;
        35: y = 16'b0011111101000010;
        36: y = 16'b0011111110011001;
        37: y = 16'b0011111111010110;
        38: y = 16'b0011111111110111;
        39: y = 16'b0011111111111110;
        40: y = 16'b0011111111101010;
        41: y = 16'b0011111110111011;
        42: y = 16'b0011111101110001;
        43: y = 16'b0011111100001100;
        44: y = 16'b0011111010001101;
        45: y = 16'b0011110111110100;
        46: y = 16'b0011110101000001;
        47: y = 16'b0011110001110011;
        48: y = 16'b0011101110001101;
        49: y = 16'b0011101010001101;
        50: y = 16'b0011100101110101;
        51: y = 16'b0011100001000100;
        52: y = 16'b0011011011111100;
        53: y = 16'b0011010110011101;
        54: y = 16'b0011010000100111;
        55: y = 16'b0011001010011011;
        56: y = 16'b0011000011111010;
        57: y = 16'b0010111101000101;
        58: y = 16'b0010110101111011;
        59: y = 16'b0010101110011110;
        60: y = 16'b0010100110101111;
        61: y = 16'b0010011110101111;
        62: y = 16'b0010010110011110;
        63: y = 16'b0010001101111101;
        64: y = 16'b0010000101001101;
        65: y = 16'b0001111100001111;
        66: y = 16'b0001110011000100;
        67: y = 16'b0001101001101101;
        68: y = 16'b0001100000001010;
        69: y = 16'b0001010110011110;
        70: y = 16'b0001001100101000;
        71: y = 16'b0001000010101011;
        72: y = 16'b0000111000100110;
        73: y = 16'b0000101110011100;
        74: y = 16'b0000100100001101;
        75: y = 16'b0000011001111001;
        76: y = 16'b0000001111100100;
        77: y = 16'b0000000101001100;
        78: y = 16'b1111111010110100;
        79: y = 16'b1111110000011100;
        80: y = 16'b1111100110000111;
        81: y = 16'b1111011011110011;
        82: y = 16'b1111010001100100;
        83: y = 16'b1111000111011010;
        84: y = 16'b1110111101010101;
        85: y = 16'b1110110011011000;
        86: y = 16'b1110101001100010;
        87: y = 16'b1110011111110110;
        88: y = 16'b1110010110010011;
        89: y = 16'b1110001100111100;
        90: y = 16'b1110000011110001;
        91: y = 16'b1101111010110011;
        92: y = 16'b1101110010000011;
        93: y = 16'b1101101001100010;
        94: y = 16'b1101100001010001;
        95: y = 16'b1101011001010001;
        96: y = 16'b1101010001100010;
        97: y = 16'b1101001010000101;
        98: y = 16'b1101000010111011;
        99: y = 16'b1100111100000110;
        100: y = 16'b1100110101100101;
        101: y = 16'b1100101111011001;
        102: y = 16'b1100101001100011;
        103: y = 16'b1100100100000100;
        104: y = 16'b1100011110111100;
        105: y = 16'b1100011010001011;
        106: y = 16'b1100010101110011;
        107: y = 16'b1100010001110011;
        108: y = 16'b1100001110001101;
        109: y = 16'b1100001010111111;
        110: y = 16'b1100001000001100;
        111: y = 16'b1100000101110011;
        112: y = 16'b1100000011110100;
        113: y = 16'b1100000010001111;
        114: y = 16'b1100000001000101;
        115: y = 16'b1100000000010110;
        116: y = 16'b1100000000000010;
        117: y = 16'b1100000000001001;
        118: y = 16'b1100000000101010;
        119: y = 16'b1100000001100111;
        120: y = 16'b1100000010111110;
        121: y = 16'b1100000100110000;
        122: y = 16'b1100000110111100;
        123: y = 16'b1100001001100010;
        124: y = 16'b1100001100100011;
        125: y = 16'b1100001111111101;
        126: y = 16'b1100010011110000;
        127: y = 16'b1100010111111100;
        128: y = 16'b1100011100100001;
        129: y = 16'b1100100001011101;
        130: y = 16'b1100100110110001;
        131: y = 16'b1100101100011011;
        132: y = 16'b1100110010011100;
        133: y = 16'b1100111000110011;
        134: y = 16'b1100111111011110;
        135: y = 16'b1101000110011110;
        136: y = 16'b1101001101110001;
        137: y = 16'b1101010101010111;
        138: y = 16'b1101011101001111;
        139: y = 16'b1101100101011000;
        140: y = 16'b1101101101110001;
        141: y = 16'b1101110110011010;
        142: y = 16'b1101111111010001;
        143: y = 16'b1110001000010101;
        144: y = 16'b1110010001100110;
        145: y = 16'b1110011011000011;
        146: y = 16'b1110100100101011;
        147: y = 16'b1110101110011100;
        148: y = 16'b1110111000010101;
        149: y = 16'b1111000010010110;
        150: y = 16'b1111001100011110;
        151: y = 16'b1111010110101011;
        152: y = 16'b1111100000111101;
        153: y = 16'b1111101011010001;
        154: y = 16'b1111110101101000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=440.0Hz, Fs=64453Hz, 16-bit

module lut_A
(
    input        [ 7:0] x,
    output       [ 7:0] x_max,
    output logic [15:0] y
);

    assign x_max = 145;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001011000001;
        2: y = 16'b0000010110000000;
        3: y = 16'b0000100000111101;
        4: y = 16'b0000101011110110;
        5: y = 16'b0000110110101010;
        6: y = 16'b0001000001010111;
        7: y = 16'b0001001011111101;
        8: y = 16'b0001010110011010;
        9: y = 16'b0001100000101100;
        10: y = 16'b0001101010110011;
        11: y = 16'b0001110100101101;
        12: y = 16'b0001111110011010;
        13: y = 16'b0010000111110111;
        14: y = 16'b0010010001000100;
        15: y = 16'b0010011010000000;
        16: y = 16'b0010100010101010;
        17: y = 16'b0010101011000001;
        18: y = 16'b0010110011000011;
        19: y = 16'b0010111010110000;
        20: y = 16'b0011000010000111;
        21: y = 16'b0011001001000111;
        22: y = 16'b0011001111101111;
        23: y = 16'b0011010101111111;
        24: y = 16'b0011011011110101;
        25: y = 16'b0011100001010001;
        26: y = 16'b0011100110010011;
        27: y = 16'b0011101010111001;
        28: y = 16'b0011101111000011;
        29: y = 16'b0011110010110001;
        30: y = 16'b0011110110000010;
        31: y = 16'b0011111000110110;
        32: y = 16'b0011111011001101;
        33: y = 16'b0011111101000110;
        34: y = 16'b0011111110100000;
        35: y = 16'b0011111111011101;
        36: y = 16'b0011111111111011;
        37: y = 16'b0011111111111011;
        38: y = 16'b0011111111011101;
        39: y = 16'b0011111110100000;
        40: y = 16'b0011111101000110;
        41: y = 16'b0011111011001101;
        42: y = 16'b0011111000110110;
        43: y = 16'b0011110110000010;
        44: y = 16'b0011110010110001;
        45: y = 16'b0011101111000011;
        46: y = 16'b0011101010111001;
        47: y = 16'b0011100110010011;
        48: y = 16'b0011100001010001;
        49: y = 16'b0011011011110101;
        50: y = 16'b0011010101111111;
        51: y = 16'b0011001111101111;
        52: y = 16'b0011001001000111;
        53: y = 16'b0011000010000111;
        54: y = 16'b0010111010110000;
        55: y = 16'b0010110011000011;
        56: y = 16'b0010101011000001;
        57: y = 16'b0010100010101010;
        58: y = 16'b0010011010000000;
        59: y = 16'b0010010001000100;
        60: y = 16'b0010000111110111;
        61: y = 16'b0001111110011010;
        62: y = 16'b0001110100101101;
        63: y = 16'b0001101010110011;
        64: y = 16'b0001100000101100;
        65: y = 16'b0001010110011010;
        66: y = 16'b0001001011111101;
        67: y = 16'b0001000001010111;
        68: y = 16'b0000110110101010;
        69: y = 16'b0000101011110110;
        70: y = 16'b0000100000111101;
        71: y = 16'b0000010110000000;
        72: y = 16'b0000001011000001;
        73: y = 16'b0000000000000000;
        74: y = 16'b1111110100111111;
        75: y = 16'b1111101010000000;
        76: y = 16'b1111011111000011;
        77: y = 16'b1111010100001010;
        78: y = 16'b1111001001010110;
        79: y = 16'b1110111110101001;
        80: y = 16'b1110110100000011;
        81: y = 16'b1110101001100110;
        82: y = 16'b1110011111010100;
        83: y = 16'b1110010101001101;
        84: y = 16'b1110001011010011;
        85: y = 16'b1110000001100110;
        86: y = 16'b1101111000001001;
        87: y = 16'b1101101110111100;
        88: y = 16'b1101100110000000;
        89: y = 16'b1101011101010110;
        90: y = 16'b1101010100111111;
        91: y = 16'b1101001100111101;
        92: y = 16'b1101000101010000;
        93: y = 16'b1100111101111001;
        94: y = 16'b1100110110111001;
        95: y = 16'b1100110000010001;
        96: y = 16'b1100101010000001;
        97: y = 16'b1100100100001011;
        98: y = 16'b1100011110101111;
        99: y = 16'b1100011001101101;
        100: y = 16'b1100010101000111;
        101: y = 16'b1100010000111101;
        102: y = 16'b1100001101001111;
        103: y = 16'b1100001001111110;
        104: y = 16'b1100000111001010;
        105: y = 16'b1100000100110011;
        106: y = 16'b1100000010111010;
        107: y = 16'b1100000001100000;
        108: y = 16'b1100000000100011;
        109: y = 16'b1100000000000101;
        110: y = 16'b1100000000000101;
        111: y = 16'b1100000000100011;
        112: y = 16'b1100000001100000;
        113: y = 16'b1100000010111010;
        114: y = 16'b1100000100110011;
        115: y = 16'b1100000111001010;
        116: y = 16'b1100001001111110;
        117: y = 16'b1100001101001111;
        118: y = 16'b1100010000111101;
        119: y = 16'b1100010101000111;
        120: y = 16'b1100011001101101;
        121: y = 16'b1100011110101111;
        122: y = 16'b1100100100001011;
        123: y = 16'b1100101010000001;
        124: y = 16'b1100110000010001;
        125: y = 16'b1100110110111001;
        126: y = 16'b1100111101111001;
        127: y = 16'b1101000101010000;
        128: y = 16'b1101001100111101;
        129: y = 16'b1101010100111111;
        130: y = 16'b1101011101010110;
        131: y = 16'b1101100110000000;
        132: y = 16'b1101101110111100;
        133: y = 16'b1101111000001001;
        134: y = 16'b1110000001100110;
        135: y = 16'b1110001011010011;
        136: y = 16'b1110010101001101;
        137: y = 16'b1110011111010100;
        138: y = 16'b1110101001100110;
        139: y = 16'b1110110100000011;
        140: y = 16'b1110111110101001;
        141: y = 16'b1111001001010110;
        142: y = 16'b1111010100001010;
        143: y = 16'b1111011111000011;
        144: y = 16'b1111101010000000;
        145: y = 16'b1111110100111111;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=466.16Hz, Fs=64453Hz, 16-bit

module lut_As
(
    input        [ 7:0] x,
    output       [ 7:0] x_max,
    output logic [15:0] y
);

    assign x_max = 137;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001011101010;
        2: y = 16'b0000010111010010;
        3: y = 16'b0000100010110111;
        4: y = 16'b0000101110010111;
        5: y = 16'b0000111001110001;
        6: y = 16'b0001000101000100;
        7: y = 16'b0001010000001110;
        8: y = 16'b0001011011001100;
        9: y = 16'b0001100101111111;
        10: y = 16'b0001110000100100;
        11: y = 16'b0001111010111010;
        12: y = 16'b0010000101000000;
        13: y = 16'b0010001110110101;
        14: y = 16'b0010011000010110;
        15: y = 16'b0010100001100011;
        16: y = 16'b0010101010011011;
        17: y = 16'b0010110010111100;
        18: y = 16'b0010111011000101;
        19: y = 16'b0011000010110110;
        20: y = 16'b0011001010001101;
        21: y = 16'b0011010001001000;
        22: y = 16'b0011010111101001;
        23: y = 16'b0011011101101100;
        24: y = 16'b0011100011010010;
        25: y = 16'b0011101000011010;
        26: y = 16'b0011101101000011;
        27: y = 16'b0011110001001101;
        28: y = 16'b0011110100110111;
        29: y = 16'b0011111000000000;
        30: y = 16'b0011111010101000;
        31: y = 16'b0011111100101111;
        32: y = 16'b0011111110010101;
        33: y = 16'b0011111111011001;
        34: y = 16'b0011111111111011;
        35: y = 16'b0011111111111011;
        36: y = 16'b0011111111011001;
        37: y = 16'b0011111110010101;
        38: y = 16'b0011111100101111;
        39: y = 16'b0011111010101000;
        40: y = 16'b0011111000000000;
        41: y = 16'b0011110100110111;
        42: y = 16'b0011110001001101;
        43: y = 16'b0011101101000011;
        44: y = 16'b0011101000011010;
        45: y = 16'b0011100011010010;
        46: y = 16'b0011011101101100;
        47: y = 16'b0011010111101001;
        48: y = 16'b0011010001001000;
        49: y = 16'b0011001010001101;
        50: y = 16'b0011000010110110;
        51: y = 16'b0010111011000101;
        52: y = 16'b0010110010111100;
        53: y = 16'b0010101010011011;
        54: y = 16'b0010100001100011;
        55: y = 16'b0010011000010110;
        56: y = 16'b0010001110110101;
        57: y = 16'b0010000101000000;
        58: y = 16'b0001111010111010;
        59: y = 16'b0001110000100100;
        60: y = 16'b0001100101111111;
        61: y = 16'b0001011011001100;
        62: y = 16'b0001010000001110;
        63: y = 16'b0001000101000100;
        64: y = 16'b0000111001110001;
        65: y = 16'b0000101110010111;
        66: y = 16'b0000100010110111;
        67: y = 16'b0000010111010010;
        68: y = 16'b0000001011101010;
        69: y = 16'b0000000000000000;
        70: y = 16'b1111110100010110;
        71: y = 16'b1111101000101110;
        72: y = 16'b1111011101001001;
        73: y = 16'b1111010001101001;
        74: y = 16'b1111000110001111;
        75: y = 16'b1110111010111100;
        76: y = 16'b1110101111110010;
        77: y = 16'b1110100100110100;
        78: y = 16'b1110011010000001;
        79: y = 16'b1110001111011100;
        80: y = 16'b1110000101000110;
        81: y = 16'b1101111011000000;
        82: y = 16'b1101110001001011;
        83: y = 16'b1101100111101010;
        84: y = 16'b1101011110011101;
        85: y = 16'b1101010101100101;
        86: y = 16'b1101001101000100;
        87: y = 16'b1101000100111011;
        88: y = 16'b1100111101001010;
        89: y = 16'b1100110101110011;
        90: y = 16'b1100101110111000;
        91: y = 16'b1100101000010111;
        92: y = 16'b1100100010010100;
        93: y = 16'b1100011100101110;
        94: y = 16'b1100010111100110;
        95: y = 16'b1100010010111101;
        96: y = 16'b1100001110110011;
        97: y = 16'b1100001011001001;
        98: y = 16'b1100001000000000;
        99: y = 16'b1100000101011000;
        100: y = 16'b1100000011010001;
        101: y = 16'b1100000001101011;
        102: y = 16'b1100000000100111;
        103: y = 16'b1100000000000101;
        104: y = 16'b1100000000000101;
        105: y = 16'b1100000000100111;
        106: y = 16'b1100000001101011;
        107: y = 16'b1100000011010001;
        108: y = 16'b1100000101011000;
        109: y = 16'b1100001000000000;
        110: y = 16'b1100001011001001;
        111: y = 16'b1100001110110011;
        112: y = 16'b1100010010111101;
        113: y = 16'b1100010111100110;
        114: y = 16'b1100011100101110;
        115: y = 16'b1100100010010100;
        116: y = 16'b1100101000010111;
        117: y = 16'b1100101110111000;
        118: y = 16'b1100110101110011;
        119: y = 16'b1100111101001010;
        120: y = 16'b1101000100111011;
        121: y = 16'b1101001101000100;
        122: y = 16'b1101010101100101;
        123: y = 16'b1101011110011101;
        124: y = 16'b1101100111101010;
        125: y = 16'b1101110001001011;
        126: y = 16'b1101111011000000;
        127: y = 16'b1110000101000110;
        128: y = 16'b1110001111011100;
        129: y = 16'b1110011010000001;
        130: y = 16'b1110100100110100;
        131: y = 16'b1110101111110010;
        132: y = 16'b1110111010111100;
        133: y = 16'b1111000110001111;
        134: y = 16'b1111010001101001;
        135: y = 16'b1111011101001001;
        136: y = 16'b1111101000101110;
        137: y = 16'b1111110100010110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=493.88Hz, Fs=64453Hz, 16-bit

module lut_B
(
    input        [ 7:0] x,
    output       [ 7:0] x_max,
    output logic [15:0] y
);

    assign x_max = 129;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001100011000;
        2: y = 16'b0000011000101101;
        3: y = 16'b0000100100111111;
        4: y = 16'b0000110001001100;
        5: y = 16'b0000111101010001;
        6: y = 16'b0001001001001101;
        7: y = 16'b0001010100111110;
        8: y = 16'b0001100000100010;
        9: y = 16'b0001101011111000;
        10: y = 16'b0001110110111110;
        11: y = 16'b0010000001110010;
        12: y = 16'b0010001100010010;
        13: y = 16'b0010010110011110;
        14: y = 16'b0010100000010011;
        15: y = 16'b0010101001110000;
        16: y = 16'b0010110010110100;
        17: y = 16'b0010111011011101;
        18: y = 16'b0011000011101010;
        19: y = 16'b0011001011011010;
        20: y = 16'b0011010010101011;
        21: y = 16'b0011011001011101;
        22: y = 16'b0011011111101110;
        23: y = 16'b0011100101011110;
        24: y = 16'b0011101010101100;
        25: y = 16'b0011101111010110;
        26: y = 16'b0011110011011101;
        27: y = 16'b0011110111000000;
        28: y = 16'b0011111001111101;
        29: y = 16'b0011111100010101;
        30: y = 16'b0011111110001000;
        31: y = 16'b0011111111010100;
        32: y = 16'b0011111111111010;
        33: y = 16'b0011111111111010;
        34: y = 16'b0011111111010100;
        35: y = 16'b0011111110001000;
        36: y = 16'b0011111100010101;
        37: y = 16'b0011111001111101;
        38: y = 16'b0011110111000000;
        39: y = 16'b0011110011011101;
        40: y = 16'b0011101111010110;
        41: y = 16'b0011101010101100;
        42: y = 16'b0011100101011110;
        43: y = 16'b0011011111101110;
        44: y = 16'b0011011001011101;
        45: y = 16'b0011010010101011;
        46: y = 16'b0011001011011010;
        47: y = 16'b0011000011101010;
        48: y = 16'b0010111011011101;
        49: y = 16'b0010110010110100;
        50: y = 16'b0010101001110000;
        51: y = 16'b0010100000010011;
        52: y = 16'b0010010110011110;
        53: y = 16'b0010001100010010;
        54: y = 16'b0010000001110010;
        55: y = 16'b0001110110111110;
        56: y = 16'b0001101011111000;
        57: y = 16'b0001100000100010;
        58: y = 16'b0001010100111110;
        59: y = 16'b0001001001001101;
        60: y = 16'b0000111101010001;
        61: y = 16'b0000110001001100;
        62: y = 16'b0000100100111111;
        63: y = 16'b0000011000101101;
        64: y = 16'b0000001100011000;
        65: y = 16'b0000000000000000;
        66: y = 16'b1111110011101000;
        67: y = 16'b1111100111010011;
        68: y = 16'b1111011011000001;
        69: y = 16'b1111001110110100;
        70: y = 16'b1111000010101111;
        71: y = 16'b1110110110110011;
        72: y = 16'b1110101011000010;
        73: y = 16'b1110011111011110;
        74: y = 16'b1110010100001000;
        75: y = 16'b1110001001000010;
        76: y = 16'b1101111110001110;
        77: y = 16'b1101110011101110;
        78: y = 16'b1101101001100010;
        79: y = 16'b1101011111101101;
        80: y = 16'b1101010110010000;
        81: y = 16'b1101001101001100;
        82: y = 16'b1101000100100011;
        83: y = 16'b1100111100010110;
        84: y = 16'b1100110100100110;
        85: y = 16'b1100101101010101;
        86: y = 16'b1100100110100011;
        87: y = 16'b1100100000010010;
        88: y = 16'b1100011010100010;
        89: y = 16'b1100010101010100;
        90: y = 16'b1100010000101010;
        91: y = 16'b1100001100100011;
        92: y = 16'b1100001001000000;
        93: y = 16'b1100000110000011;
        94: y = 16'b1100000011101011;
        95: y = 16'b1100000001111000;
        96: y = 16'b1100000000101100;
        97: y = 16'b1100000000000110;
        98: y = 16'b1100000000000110;
        99: y = 16'b1100000000101100;
        100: y = 16'b1100000001111000;
        101: y = 16'b1100000011101011;
        102: y = 16'b1100000110000011;
        103: y = 16'b1100001001000000;
        104: y = 16'b1100001100100011;
        105: y = 16'b1100010000101010;
        106: y = 16'b1100010101010100;
        107: y = 16'b1100011010100010;
        108: y = 16'b1100100000010010;
        109: y = 16'b1100100110100011;
        110: y = 16'b1100101101010101;
        111: y = 16'b1100110100100110;
        112: y = 16'b1100111100010110;
        113: y = 16'b1101000100100011;
        114: y = 16'b1101001101001100;
        115: y = 16'b1101010110010000;
        116: y = 16'b1101011111101101;
        117: y = 16'b1101101001100010;
        118: y = 16'b1101110011101110;
        119: y = 16'b1101111110001110;
        120: y = 16'b1110001001000010;
        121: y = 16'b1110010100001000;
        122: y = 16'b1110011111011110;
        123: y = 16'b1110101011000010;
        124: y = 16'b1110110110110011;
        125: y = 16'b1111000010101111;
        126: y = 16'b1111001110110100;
        127: y = 16'b1111011011000001;
        128: y = 16'b1111100111010011;
        129: y = 16'b1111110011101000;
        default: y = 16'b0;
        endcase

endmodule

