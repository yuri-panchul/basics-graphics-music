//Copyright (C)2014-2025 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.11.03 Education
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9
//Device Version: C
//Created Time: Wed Dec 31 16:15:04 2025

module Gowin_SDPB (dout, clka, cea, reseta, clkb, ceb, resetb, oce, ada, din, adb);

output [7:0] dout;
input clka;
input cea;
input reseta;
input clkb;
input ceb;
input resetb;
input oce;
input [12:0] ada;
input [7:0] din;
input [12:0] adb;

wire [27:0] sdpb_inst_0_dout_w;
wire [3:0] sdpb_inst_0_dout;
wire [27:0] sdpb_inst_1_dout_w;
wire [7:4] sdpb_inst_1_dout;
wire [23:0] sdpb_inst_2_dout_w;
wire [7:0] sdpb_inst_2_dout;
wire dff_q_0;
wire gw_gnd;

assign gw_gnd = 1'b0;

SDPB sdpb_inst_0 (
    .DO({sdpb_inst_0_dout_w[27:0],sdpb_inst_0_dout[3:0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[12]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[12]}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3:0]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd})
);

defparam sdpb_inst_0.READ_MODE = 1'b0;
defparam sdpb_inst_0.BIT_WIDTH_0 = 4;
defparam sdpb_inst_0.BIT_WIDTH_1 = 4;
defparam sdpb_inst_0.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_0.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_0.RESET_MODE = "SYNC";
defparam sdpb_inst_0.INIT_RAM_00 = 256'h0F404530C49C507E93390941025454353EF30C45D1049302FCF40D53090D52FC;
defparam sdpb_inst_0.INIT_RAM_01 = 256'h50450E1519C101E71D052FCF4045052F21C04504E549493E902F0D5404FD3595;
defparam sdpb_inst_0.INIT_RAM_02 = 256'hE0392F21C0F3D1CC50EF9414932585045243FE039510CD19E560D9E9D0410D9E;
defparam sdpb_inst_0.INIT_RAM_03 = 256'hE902FCF405252905451039540E415153EF30F4FDDF3015085009519C10450939;
defparam sdpb_inst_0.INIT_RAM_04 = 256'hE0419756055052FCF40D5CC9305335049C560541405CF60E9049254E58520520;
defparam sdpb_inst_0.INIT_RAM_05 = 256'h30C4E549F200EFE041414905304135133F04E9302554053850E2541921001CC5;
defparam sdpb_inst_0.INIT_RAM_06 = 256'h2FCED52F21C04350490D9E1049CCFD04E5253540193966F0951010C530E904E5;
defparam sdpb_inst_0.INIT_RAM_07 = 256'h5950F404530C49C507E93390941025454353EF30C45D1049302FCF40D53090D5;
defparam sdpb_inst_0.INIT_RAM_08 = 256'hD9E50450E1519C101E71D052FCF4045052F21C04504E549493E902F0D5404FD3;
defparam sdpb_inst_0.INIT_RAM_09 = 256'h939E0392F21C0F3D1CC50EF9414932585045243FE039510CD19E560D9E9D0410;
defparam sdpb_inst_0.INIT_RAM_0A = 256'h520E902FCF405252905451039540E415153EF30F4FDDF3015085009519C10450;
defparam sdpb_inst_0.INIT_RAM_0B = 256'hCC5E0419756055052FCF40D5CC9305335049C560541405CF60E9049254E58520;
defparam sdpb_inst_0.INIT_RAM_0C = 256'h4E530C4E549F200EFE041414905304135133F04E9302554053850E2541921001;
defparam sdpb_inst_0.INIT_RAM_0D = 256'h0D52FCED52F21C04350490D9E1049CCFD04E5253540193966F0951010C530E90;
defparam sdpb_inst_0.INIT_RAM_0E = 256'hFD35950F404530C49C507E93390941025454353EF30C45D1049302FCF40D5309;
defparam sdpb_inst_0.INIT_RAM_0F = 256'h410D9E50450E1519C101E71D052FCF4045052F21C04504E549493E902F0D5404;
defparam sdpb_inst_0.INIT_RAM_10 = 256'h450939E0392F21C0F3D1CC50EF9414932585045243FE039510CD19E560D9E9D0;
defparam sdpb_inst_0.INIT_RAM_11 = 256'h520520E902FCF405252905451039540E415153EF30F4FDDF3015085009519C10;
defparam sdpb_inst_0.INIT_RAM_12 = 256'h001CC5E0419756055052FCF40D5CC9305335049C560541405CF60E9049254E58;
defparam sdpb_inst_0.INIT_RAM_13 = 256'hE904E530C4E549F200EFE041414905304135133F04E9302554053850E2541921;
defparam sdpb_inst_0.INIT_RAM_14 = 256'h3090D52FCED52F21C04350490D9E1049CCFD04E5253540193966F0951010C530;
defparam sdpb_inst_0.INIT_RAM_15 = 256'h404FD35950F404530C49C507E93390941025454353EF30C45D1049302FCF40D5;
defparam sdpb_inst_0.INIT_RAM_16 = 256'h9D0410D9E50450E1519C101E71D052FCF4045052F21C04504E549493E902F0D5;
defparam sdpb_inst_0.INIT_RAM_17 = 256'hC10450939E0392F21C0F3D1CC50EF9414932585045243FE039510CD19E560D9E;
defparam sdpb_inst_0.INIT_RAM_18 = 256'hE58520520E902FCF405252905451039540E415153EF30F4FDDF3015085009519;
defparam sdpb_inst_0.INIT_RAM_19 = 256'h921001CC5E0419756055052FCF40D5CC9305335049C560541405CF60E9049254;
defparam sdpb_inst_0.INIT_RAM_1A = 256'h530E904E530C4E549F200EFE041414905304135133F04E9302554053850E2541;
defparam sdpb_inst_0.INIT_RAM_1B = 256'h0D53090D52FCED52F21C04350490D9E1049CCFD04E5253540193966F0951010C;
defparam sdpb_inst_0.INIT_RAM_1C = 256'h0D5404FD35950F404530C49C507E93390941025454353EF30C45D1049302FCF4;
defparam sdpb_inst_0.INIT_RAM_1D = 256'hD9E9D0410D9E50450E1519C101E71D052FCF4045052F21C04504E549493E902F;
defparam sdpb_inst_0.INIT_RAM_1E = 256'h519C10450939E0392F21C0F3D1CC50EF9414932585045243FE039510CD19E560;
defparam sdpb_inst_0.INIT_RAM_1F = 256'h254E58520520E902FCF405252905451039540E415153EF30F4FDDF3015085009;
defparam sdpb_inst_0.INIT_RAM_20 = 256'h541921001CC5E0419756055052FCF40D5CC9305335049C560541405CF60E9049;
defparam sdpb_inst_0.INIT_RAM_21 = 256'h10C530E904E530C4E549F200EFE041414905304135133F04E9302554053850E2;
defparam sdpb_inst_0.INIT_RAM_22 = 256'hCF40D53090D52FCED52F21C04350490D9E1049CCFD04E5253540193966F09510;
defparam sdpb_inst_0.INIT_RAM_23 = 256'h02F0D5404FD35950F404530C49C507E93390941025454353EF30C45D1049302F;
defparam sdpb_inst_0.INIT_RAM_24 = 256'h560D9E9D0410D9E50450E1519C101E71D052FCF4045052F21C04504E549493E9;
defparam sdpb_inst_0.INIT_RAM_25 = 256'h009519C10450939E0392F21C0F3D1CC50EF9414932585045243FE039510CD19E;
defparam sdpb_inst_0.INIT_RAM_26 = 256'h049254E58520520E902FCF405252905451039540E415153EF30F4FDDF3015085;
defparam sdpb_inst_0.INIT_RAM_27 = 256'h0E2541921001CC5E0419756055052FCF40D5CC9305335049C560541405CF60E9;
defparam sdpb_inst_0.INIT_RAM_28 = 256'h51010C530E904E530C4E549F200EFE041414905304135133F04E930255405385;
defparam sdpb_inst_0.INIT_RAM_29 = 256'h02FCF40D53090D52FCED52F21C04350490D9E1049CCFD04E5253540193966F09;
defparam sdpb_inst_0.INIT_RAM_2A = 256'h3E902F0D5404FD35950F404530C49C507E93390941025454353EF30C45D10493;
defparam sdpb_inst_0.INIT_RAM_2B = 256'h19E560D9E9D0410D9E50450E1519C101E71D052FCF4045052F21C04504E54949;
defparam sdpb_inst_0.INIT_RAM_2C = 256'h085009519C10450939E0392F21C0F3D1CC50EF9414932585045243FE039510CD;
defparam sdpb_inst_0.INIT_RAM_2D = 256'h0E9049254E58520520E902FCF405252905451039540E415153EF30F4FDDF3015;
defparam sdpb_inst_0.INIT_RAM_2E = 256'h3850E2541921001CC5E0419756055052FCF40D5CC9305335049C560541405CF6;
defparam sdpb_inst_0.INIT_RAM_2F = 256'hF0951010C530E904E530C4E549F200EFE041414905304135133F04E930255405;
defparam sdpb_inst_0.INIT_RAM_30 = 256'h49302FCF40D53090D52FCED52F21C04350490D9E1049CCFD04E5253540193966;
defparam sdpb_inst_0.INIT_RAM_31 = 256'h9493E902F0D5404FD35950F404530C49C507E93390941025454353EF30C45D10;
defparam sdpb_inst_0.INIT_RAM_32 = 256'h0CD19E560D9E9D0410D9E50450E1519C101E71D052FCF4045052F21C04504E54;
defparam sdpb_inst_0.INIT_RAM_33 = 256'h015085009519C10450939E0392F21C0F3D1CC50EF9414932585045243FE03951;
defparam sdpb_inst_0.INIT_RAM_34 = 256'hCF60E9049254E58520520E902FCF405252905451039540E415153EF30F4FDDF3;
defparam sdpb_inst_0.INIT_RAM_35 = 256'h4053850E2541921001CC5E0419756055052FCF40D5CC9305335049C560541405;
defparam sdpb_inst_0.INIT_RAM_36 = 256'h966F0951010C530E904E530C4E549F200EFE041414905304135133F04E930255;
defparam sdpb_inst_0.INIT_RAM_37 = 256'hD1049302FCF40D53090D52FCED52F21C04350490D9E1049CCFD04E5253540193;
defparam sdpb_inst_0.INIT_RAM_38 = 256'hE549493E902F0D5404FD35950F404530C49C507E93390941025454353EF30C45;
defparam sdpb_inst_0.INIT_RAM_39 = 256'h9510CD19E560D9E9D0410D9E50450E1519C101E71D052FCF4045052F21C04504;
defparam sdpb_inst_0.INIT_RAM_3A = 256'hDF3015085009519C10450939E0392F21C0F3D1CC50EF9414932585045243FE03;
defparam sdpb_inst_0.INIT_RAM_3B = 256'h405CF60E9049254E58520520E902FCF405252905451039540E415153EF30F4FD;
defparam sdpb_inst_0.INIT_RAM_3C = 256'h2554053850E2541921001CC5E0419756055052FCF40D5CC9305335049C560541;
defparam sdpb_inst_0.INIT_RAM_3D = 256'h193966F0951010C530E904E530C4E549F200EFE041414905304135133F04E930;
defparam sdpb_inst_0.INIT_RAM_3E = 256'hC45D1049302FCF40D53090D52FCED52F21C04350490D9E1049CCFD04E5253540;
defparam sdpb_inst_0.INIT_RAM_3F = 256'h504E549493E902F0D5404FD35950F404530C49C507E93390941025454353EF30;

SDPB sdpb_inst_1 (
    .DO({sdpb_inst_1_dout_w[27:0],sdpb_inst_1_dout[7:4]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[12]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[12]}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:4]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd})
);

defparam sdpb_inst_1.READ_MODE = 1'b0;
defparam sdpb_inst_1.BIT_WIDTH_0 = 4;
defparam sdpb_inst_1.BIT_WIDTH_1 = 4;
defparam sdpb_inst_1.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_1.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_1.RESET_MODE = "SYNC";
defparam sdpb_inst_1.INIT_RAM_00 = 256'h2662667227666266667676662777676676662276662767276666267776266764;
defparam sdpb_inst_1.INIT_RAM_01 = 256'h6275226776662666662676666276267666627727676666666276766726667766;
defparam sdpb_inst_1.INIT_RAM_02 = 256'h6276766662666666726667676676762677776627677226666672666662662666;
defparam sdpb_inst_1.INIT_RAM_03 = 256'h6627666626777626776276742276776766626666666266276276776662772676;
defparam sdpb_inst_1.INIT_RAM_04 = 256'h6276667627626766662676666267762766672676777667266276766666677672;
defparam sdpb_inst_1.INIT_RAM_05 = 256'h7227666667726662767666776276666666276672776776674227776676726667;
defparam sdpb_inst_1.INIT_RAM_06 = 256'h7642677666627762662666627666662767767662666666626772676762662767;
defparam sdpb_inst_1.INIT_RAM_07 = 256'h7662662667227666266667676662777676676662276662767276666267776266;
defparam sdpb_inst_1.INIT_RAM_08 = 256'h6666275226776662666662676666276267666627727676666666276766726667;
defparam sdpb_inst_1.INIT_RAM_09 = 256'h6766276766662666666726667676676762677776627677226666672666662662;
defparam sdpb_inst_1.INIT_RAM_0A = 256'h6726627666626777626776276742276776766626666666266276276776662772;
defparam sdpb_inst_1.INIT_RAM_0B = 256'h6676276667627626766662676666267762766672676777667266276766666677;
defparam sdpb_inst_1.INIT_RAM_0C = 256'h7677227666667726662767666776276666666276672776776674227776676726;
defparam sdpb_inst_1.INIT_RAM_0D = 256'h2667642677666627762662666627666662767767662666666626772676762662;
defparam sdpb_inst_1.INIT_RAM_0E = 256'h6677662662667227666266667676662777676676662276662767276666267776;
defparam sdpb_inst_1.INIT_RAM_0F = 256'h6626666275226776662666662676666276267666627727676666666276766726;
defparam sdpb_inst_1.INIT_RAM_10 = 256'h7726766276766662666666726667676676762677776627677226666672666662;
defparam sdpb_inst_1.INIT_RAM_11 = 256'h6776726627666626777626776276742276776766626666666266276276776662;
defparam sdpb_inst_1.INIT_RAM_12 = 256'h7266676276667627626766662676666267762766672676777667266276766666;
defparam sdpb_inst_1.INIT_RAM_13 = 256'h6627677227666667726662767666776276666666276672776776674227776676;
defparam sdpb_inst_1.INIT_RAM_14 = 256'h7762667642677666627762662666627666662767767662666666626772676762;
defparam sdpb_inst_1.INIT_RAM_15 = 256'h7266677662662667227666266667676662777676676662276662767276666267;
defparam sdpb_inst_1.INIT_RAM_16 = 256'h6626626666275226776662666662676666276267666627727676666666276766;
defparam sdpb_inst_1.INIT_RAM_17 = 256'h6627726766276766662666666726667676676762677776627677226666672666;
defparam sdpb_inst_1.INIT_RAM_18 = 256'h6666776726627666626777626776276742276776766626666666266276276776;
defparam sdpb_inst_1.INIT_RAM_19 = 256'h6767266676276667627626766662676666267762766672676777667266276766;
defparam sdpb_inst_1.INIT_RAM_1A = 256'h7626627677227666667726662767666776276666666276672776776674227776;
defparam sdpb_inst_1.INIT_RAM_1B = 256'h2677762667642677666627762662666627666662767767662666666626772676;
defparam sdpb_inst_1.INIT_RAM_1C = 256'h7667266677662662667227666266667676662777676676662276662767276666;
defparam sdpb_inst_1.INIT_RAM_1D = 256'h6666626626666275226776662666662676666276267666627727676666666276;
defparam sdpb_inst_1.INIT_RAM_1E = 256'h7766627726766276766662666666726667676676762677776627677226666672;
defparam sdpb_inst_1.INIT_RAM_1F = 256'h7666666776726627666626777626776276742276776766626666666266276276;
defparam sdpb_inst_1.INIT_RAM_20 = 256'h7766767266676276667627626766662676666267762766672676777667266276;
defparam sdpb_inst_1.INIT_RAM_21 = 256'h6767626627677227666667726662767666776276666666276672776776674227;
defparam sdpb_inst_1.INIT_RAM_22 = 256'h6662677762667642677666627762662666627666662767767662666666626772;
defparam sdpb_inst_1.INIT_RAM_23 = 256'h2767667266677662662667227666266667676662777676676662276662767276;
defparam sdpb_inst_1.INIT_RAM_24 = 256'h6726666626626666275226776662666662676666276267666627727676666666;
defparam sdpb_inst_1.INIT_RAM_25 = 256'h2767766627726766276766662666666726667676676762677776627677226666;
defparam sdpb_inst_1.INIT_RAM_26 = 256'h2767666666776726627666626777626776276742276776766626666666266276;
defparam sdpb_inst_1.INIT_RAM_27 = 256'h2277766767266676276667627626766662676666267762766672676777667266;
defparam sdpb_inst_1.INIT_RAM_28 = 256'h7726767626627677227666667726662767666776276666666276672776776674;
defparam sdpb_inst_1.INIT_RAM_29 = 256'h2766662677762667642677666627762662666627666662767767662666666626;
defparam sdpb_inst_1.INIT_RAM_2A = 256'h6662767667266677662662667227666266667676662777676676662276662767;
defparam sdpb_inst_1.INIT_RAM_2B = 256'h6666726666626626666275226776662666662676666276267666627727676666;
defparam sdpb_inst_1.INIT_RAM_2C = 256'h2762767766627726766276766662666666726667676676762677776627677226;
defparam sdpb_inst_1.INIT_RAM_2D = 256'h2662767666666776726627666626777626776276742276776766626666666266;
defparam sdpb_inst_1.INIT_RAM_2E = 256'h6742277766767266676276667627626766662676666267762766672676777667;
defparam sdpb_inst_1.INIT_RAM_2F = 256'h6267726767626627677227666667726662767666776276666666276672776776;
defparam sdpb_inst_1.INIT_RAM_30 = 256'h7672766662677762667642677666627762662666627666662767767662666666;
defparam sdpb_inst_1.INIT_RAM_31 = 256'h6666662767667266677662662667227666266667676662777676676662276662;
defparam sdpb_inst_1.INIT_RAM_32 = 256'h2266666726666626626666275226776662666662676666276267666627727676;
defparam sdpb_inst_1.INIT_RAM_33 = 256'h2662762767766627726766276766662666666726667676676762677776627677;
defparam sdpb_inst_1.INIT_RAM_34 = 256'h6672662767666666776726627666626777626776276742276776766626666666;
defparam sdpb_inst_1.INIT_RAM_35 = 256'h7766742277766767266676276667627626766662676666267762766672676777;
defparam sdpb_inst_1.INIT_RAM_36 = 256'h6666267726767626627677227666667726662767666776276666666276672776;
defparam sdpb_inst_1.INIT_RAM_37 = 256'h6627672766662677762667642677666627762662666627666662767767662666;
defparam sdpb_inst_1.INIT_RAM_38 = 256'h6766666662767667266677662662667227666266667676662777676676662276;
defparam sdpb_inst_1.INIT_RAM_39 = 256'h6772266666726666626626666275226776662666662676666276267666627727;
defparam sdpb_inst_1.INIT_RAM_3A = 256'h6662662762767766627726766276766662666666726667676676762677776627;
defparam sdpb_inst_1.INIT_RAM_3B = 256'h7776672662767666666776726627666626777626776276742276776766626666;
defparam sdpb_inst_1.INIT_RAM_3C = 256'h7767766742277766767266676276667627626766662676666267762766672676;
defparam sdpb_inst_1.INIT_RAM_3D = 256'h6666666267726767626627677227666667726662767666776276666666276672;
defparam sdpb_inst_1.INIT_RAM_3E = 256'h2766627672766662677762667642677666627762662666627666662767767662;
defparam sdpb_inst_1.INIT_RAM_3F = 256'h7276766666662767667266677662662667227666266667676662777676676662;

SDPB sdpb_inst_2 (
    .DO({sdpb_inst_2_dout_w[23:0],sdpb_inst_2_dout[7:0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,ada[12],ada[11]}),
    .BLKSELB({gw_gnd,adb[12],adb[11]}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_2.READ_MODE = 1'b0;
defparam sdpb_inst_2.BIT_WIDTH_0 = 8;
defparam sdpb_inst_2.BIT_WIDTH_1 = 8;
defparam sdpb_inst_2.BLK_SEL_0 = 3'b010;
defparam sdpb_inst_2.BLK_SEL_1 = 3'b010;
defparam sdpb_inst_2.RESET_MODE = "SYNC";
defparam sdpb_inst_2.INIT_RAM_00 = 256'h2E617571696C6120616E67616D2065726F6C6F642074652065726F62616C2074;
defparam sdpb_inst_2.INIT_RAM_01 = 256'h6E2073697571202C6D61696E6576206D696E696D206461206D696E6520745520;
defparam sdpb_inst_2.INIT_RAM_02 = 256'h6F62616C206F636D616C6C75206E6F697461746963726578652064757274736F;
defparam sdpb_inst_2.INIT_RAM_03 = 256'h646F6D6D6F632061652078652070697571696C61207475206973696E20736972;
defparam sdpb_inst_2.INIT_RAM_04 = 256'h6C6F6420657275726920657475612073697544202E7461757165736E6F63206F;
defparam sdpb_inst_2.INIT_RAM_05 = 256'h6574617470756C6F76206E692074697265646E65686572706572206E6920726F;
defparam sdpb_inst_2.INIT_RAM_06 = 256'h6775662075652065726F6C6F64206D756C6C696320657373652074696C657620;
defparam sdpb_inst_2.INIT_RAM_07 = 256'h697320727565747065637845202E727574616972617020616C6C756E20746169;
defparam sdpb_inst_2.INIT_RAM_08 = 256'h6564696F7270206E6F6E2074617461646970756320746163656163636F20746E;
defparam sdpb_inst_2.INIT_RAM_09 = 256'h6564206169636966666F206975712061706C7563206E6920746E7573202C746E;
defparam sdpb_inst_2.INIT_RAM_0A = 256'h75726F62616C20747365206469206D696E612074696C6C6F6D20746E75726573;
defparam sdpb_inst_2.INIT_RAM_0B = 256'h6F63202C74656D612074697320726F6C6F64206D75737069206D65726F4C2E6D;
defparam sdpb_inst_2.INIT_RAM_0C = 256'h6420646573202C74696C6520676E69637369706964612072757465746365736E;
defparam sdpb_inst_2.INIT_RAM_0D = 256'h6C20747520746E7564696469636E6920726F706D657420646F6D73756965206F;
defparam sdpb_inst_2.INIT_RAM_0E = 256'h7455202E617571696C6120616E67616D2065726F6C6F642074652065726F6261;
defparam sdpb_inst_2.INIT_RAM_0F = 256'h74736F6E2073697571202C6D61696E6576206D696E696D206461206D696E6520;
defparam sdpb_inst_2.INIT_RAM_10 = 256'h7369726F62616C206F636D616C6C75206E6F6974617469637265786520647572;
defparam sdpb_inst_2.INIT_RAM_11 = 256'h63206F646F6D6D6F632061652078652070697571696C61207475206973696E20;
defparam sdpb_inst_2.INIT_RAM_12 = 256'h20726F6C6F6420657275726920657475612073697544202E7461757165736E6F;
defparam sdpb_inst_2.INIT_RAM_13 = 256'h6576206574617470756C6F76206E692074697265646E65686572706572206E69;
defparam sdpb_inst_2.INIT_RAM_14 = 256'h7461696775662075652065726F6C6F64206D756C6C696320657373652074696C;
defparam sdpb_inst_2.INIT_RAM_15 = 256'h20746E697320727565747065637845202E727574616972617020616C6C756E20;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(adb[12]),
  .CLK(clkb),
  .CE(ceb)
);
MUX2 mux_inst_2 (
  .O(dout[0]),
  .I0(sdpb_inst_0_dout[0]),
  .I1(sdpb_inst_2_dout[0]),
  .S0(dff_q_0)
);
MUX2 mux_inst_5 (
  .O(dout[1]),
  .I0(sdpb_inst_0_dout[1]),
  .I1(sdpb_inst_2_dout[1]),
  .S0(dff_q_0)
);
MUX2 mux_inst_8 (
  .O(dout[2]),
  .I0(sdpb_inst_0_dout[2]),
  .I1(sdpb_inst_2_dout[2]),
  .S0(dff_q_0)
);
MUX2 mux_inst_11 (
  .O(dout[3]),
  .I0(sdpb_inst_0_dout[3]),
  .I1(sdpb_inst_2_dout[3]),
  .S0(dff_q_0)
);
MUX2 mux_inst_14 (
  .O(dout[4]),
  .I0(sdpb_inst_1_dout[4]),
  .I1(sdpb_inst_2_dout[4]),
  .S0(dff_q_0)
);
MUX2 mux_inst_17 (
  .O(dout[5]),
  .I0(sdpb_inst_1_dout[5]),
  .I1(sdpb_inst_2_dout[5]),
  .S0(dff_q_0)
);
MUX2 mux_inst_20 (
  .O(dout[6]),
  .I0(sdpb_inst_1_dout[6]),
  .I1(sdpb_inst_2_dout[6]),
  .S0(dff_q_0)
);
MUX2 mux_inst_23 (
  .O(dout[7]),
  .I0(sdpb_inst_1_dout[7]),
  .I1(sdpb_inst_2_dout[7]),
  .S0(dff_q_0)
);
endmodule //Gowin_SDPB
