`include "config.svh"

module top
# (
  parameter clk_mhz = 50,
            w_key   = 4,
            w_sw    = 8,
            w_led   = 8,
            w_digit = 8,
            w_gpio  = 20
)
(
  input                        clk,
  input                        rst,

  // Keys, switches, LEDs

  input        [w_key   - 1:0] key,
  input        [w_sw    - 1:0] sw,
  output logic [w_led   - 1:0] led,

  // A dynamic seven-segment display

  output logic [          7:0] abcdefgh,
  output logic [w_digit - 1:0] digit,

  // VGA

  output logic                 vsync,
  output logic                 hsync,
  output logic [          3:0] red,
  output logic [          3:0] green,
  output logic [          3:0] blue,

  // General-purpose Input/Output

  inout  logic [w_gpio  - 1:0] gpio
);

  //--------------------------------------------------------------------------

  // assign led      = '0;
  // assign abcdefgh = '0;
  // assign digit    = '0;
     assign vsync    = '0;
     assign hsync    = '0;
     assign red      = '0;
     assign green    = '0;
     assign blue     = '0;

  //--------------------------------------------------------------------------

  logic [31:0] cnt;

  always_ff @ (posedge clk or posedge rst)
    if (rst)
      cnt <= '0;
    else
      cnt <= cnt + 1'd1;

  wire enable = (cnt [22:0] == '0);

  //--------------------------------------------------------------------------

  wire button_on = | key;

  logic [w_led - 1:0] shift_reg;

  always_ff @ (posedge clk or posedge rst)
    if (rst)
      shift_reg <= '1;
    else if (enable)
      shift_reg <= { button_on, shift_reg [w_led - 1:1] };

  assign led      = w_led'   (shift_reg);
  assign abcdefgh = 8'       (shift_reg);
  assign digit    = w_digit' (shift_reg);

  // Exercise 1: Make the light move in the opposite direction.

  // Exercise 2: Make the light moving in a loop.
  // Use another key to reset the moving lights back to no lights.

  // Exercise 3: Display the state of the shift register
  // on a seven-segment display, moving the light in a circle.

endmodule
