// y(t) = sin(pi*F*t/2), F=261.63Hz, Fs=48828Hz, 16-bit

module table_48828_C
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 46;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001000100011;
        2: y = 16'b0000010001000110;
        3: y = 16'b0000011001101000;
        4: y = 16'b0000100010001000;
        5: y = 16'b0000101010100101;
        6: y = 16'b0000110010111111;
        7: y = 16'b0000111011010110;
        8: y = 16'b0001000011101000;
        9: y = 16'b0001001011110110;
        10: y = 16'b0001010011111110;
        11: y = 16'b0001011100000000;
        12: y = 16'b0001100011111100;
        13: y = 16'b0001101011110000;
        14: y = 16'b0001110011011101;
        15: y = 16'b0001111011000001;
        16: y = 16'b0010000010011101;
        17: y = 16'b0010001001101111;
        18: y = 16'b0010010000111000;
        19: y = 16'b0010010111110110;
        20: y = 16'b0010011110101001;
        21: y = 16'b0010100101010001;
        22: y = 16'b0010101011101101;
        23: y = 16'b0010110001111101;
        24: y = 16'b0010111000000000;
        25: y = 16'b0010111101110110;
        26: y = 16'b0011000011011111;
        27: y = 16'b0011001000111001;
        28: y = 16'b0011001110000101;
        29: y = 16'b0011010011000011;
        30: y = 16'b0011010111110001;
        31: y = 16'b0011011100010000;
        32: y = 16'b0011100000011111;
        33: y = 16'b0011100100011110;
        34: y = 16'b0011101000001101;
        35: y = 16'b0011101011101011;
        36: y = 16'b0011101110111000;
        37: y = 16'b0011110001110101;
        38: y = 16'b0011110100011111;
        39: y = 16'b0011110110111001;
        40: y = 16'b0011111001000001;
        41: y = 16'b0011111010110111;
        42: y = 16'b0011111100011011;
        43: y = 16'b0011111101101101;
        44: y = 16'b0011111110101101;
        45: y = 16'b0011111111011010;
        46: y = 16'b0011111111110110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(pi*F*t/2), F=277.18Hz, Fs=48828Hz, 16-bit

module table_48828_Cs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 44;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001000111100;
        2: y = 16'b0000010001110111;
        3: y = 16'b0000011010110000;
        4: y = 16'b0000100011101000;
        5: y = 16'b0000101100011101;
        6: y = 16'b0000110101001110;
        7: y = 16'b0000111101111011;
        8: y = 16'b0001000110100100;
        9: y = 16'b0001001111000111;
        10: y = 16'b0001010111100011;
        11: y = 16'b0001011111111001;
        12: y = 16'b0001101000001000;
        13: y = 16'b0001110000001110;
        14: y = 16'b0001111000001011;
        15: y = 16'b0001111111111111;
        16: y = 16'b0010000111101010;
        17: y = 16'b0010001111001001;
        18: y = 16'b0010010110011110;
        19: y = 16'b0010011101100110;
        20: y = 16'b0010100100100011;
        21: y = 16'b0010101011010010;
        22: y = 16'b0010110001110101;
        23: y = 16'b0010111000001001;
        24: y = 16'b0010111110001111;
        25: y = 16'b0011000100000110;
        26: y = 16'b0011001001101110;
        27: y = 16'b0011001111000110;
        28: y = 16'b0011010100001110;
        29: y = 16'b0011011001000110;
        30: y = 16'b0011011101101100;
        31: y = 16'b0011100010000001;
        32: y = 16'b0011100110000101;
        33: y = 16'b0011101001110111;
        34: y = 16'b0011101101010110;
        35: y = 16'b0011110000100011;
        36: y = 16'b0011110011011101;
        37: y = 16'b0011110110000100;
        38: y = 16'b0011111000011000;
        39: y = 16'b0011111010011001;
        40: y = 16'b0011111100000110;
        41: y = 16'b0011111101100000;
        42: y = 16'b0011111110100101;
        43: y = 16'b0011111111010111;
        44: y = 16'b0011111111110101;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(pi*F*t/2), F=293.66Hz, Fs=48828Hz, 16-bit

module table_48828_D
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 41;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001001100101;
        2: y = 16'b0000010011001000;
        3: y = 16'b0000011100101010;
        4: y = 16'b0000100110001010;
        5: y = 16'b0000101111100110;
        6: y = 16'b0000111000111110;
        7: y = 16'b0001000010010000;
        8: y = 16'b0001001011011101;
        9: y = 16'b0001010100100011;
        10: y = 16'b0001011101100001;
        11: y = 16'b0001100110010111;
        12: y = 16'b0001101111000100;
        13: y = 16'b0001110111100111;
        14: y = 16'b0001111111111111;
        15: y = 16'b0010001000001100;
        16: y = 16'b0010010000001101;
        17: y = 16'b0010011000000001;
        18: y = 16'b0010011111100111;
        19: y = 16'b0010100110111110;
        20: y = 16'b0010101110000111;
        21: y = 16'b0010110101000001;
        22: y = 16'b0010111011101010;
        23: y = 16'b0011000010000010;
        24: y = 16'b0011001000001001;
        25: y = 16'b0011001101111110;
        26: y = 16'b0011010011100000;
        27: y = 16'b0011011000110000;
        28: y = 16'b0011011101101100;
        29: y = 16'b0011100010010100;
        30: y = 16'b0011100110101001;
        31: y = 16'b0011101010101000;
        32: y = 16'b0011101110010011;
        33: y = 16'b0011110001101000;
        34: y = 16'b0011110100100111;
        35: y = 16'b0011110111010001;
        36: y = 16'b0011111001100100;
        37: y = 16'b0011111011100001;
        38: y = 16'b0011111101001000;
        39: y = 16'b0011111110011000;
        40: y = 16'b0011111111010001;
        41: y = 16'b0011111111110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(pi*F*t/2), F=311.13Hz, Fs=48828Hz, 16-bit

module table_48828_Ds
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 39;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001010000011;
        2: y = 16'b0000010100000101;
        3: y = 16'b0000011110000110;
        4: y = 16'b0000101000000011;
        5: y = 16'b0000110001111100;
        6: y = 16'b0000111011110001;
        7: y = 16'b0001000101011111;
        8: y = 16'b0001001111000111;
        9: y = 16'b0001011000100110;
        10: y = 16'b0001100001111110;
        11: y = 16'b0001101011001011;
        12: y = 16'b0001110100001110;
        13: y = 16'b0001111101000101;
        14: y = 16'b0010000101110000;
        15: y = 16'b0010001110001110;
        16: y = 16'b0010010110011110;
        17: y = 16'b0010011110011111;
        18: y = 16'b0010100110010000;
        19: y = 16'b0010101101110001;
        20: y = 16'b0010110101000001;
        21: y = 16'b0010111011111110;
        22: y = 16'b0011000010101010;
        23: y = 16'b0011001001000010;
        24: y = 16'b0011001111000110;
        25: y = 16'b0011010100110110;
        26: y = 16'b0011011010010001;
        27: y = 16'b0011011111010110;
        28: y = 16'b0011100100000101;
        29: y = 16'b0011101000011110;
        30: y = 16'b0011101100100000;
        31: y = 16'b0011110000001010;
        32: y = 16'b0011110011011101;
        33: y = 16'b0011110110011000;
        34: y = 16'b0011111000111010;
        35: y = 16'b0011111011000100;
        36: y = 16'b0011111100110101;
        37: y = 16'b0011111110001101;
        38: y = 16'b0011111111001100;
        39: y = 16'b0011111111110010;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(pi*F*t/2), F=329.63Hz, Fs=48828Hz, 16-bit

module table_48828_E
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 37;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001010100101;
        2: y = 16'b0000010101001001;
        3: y = 16'b0000011111101010;
        4: y = 16'b0000101010001001;
        5: y = 16'b0000110100100010;
        6: y = 16'b0000111110110110;
        7: y = 16'b0001001001000011;
        8: y = 16'b0001010011001000;
        9: y = 16'b0001011101000011;
        10: y = 16'b0001100110110101;
        11: y = 16'b0001110000011011;
        12: y = 16'b0001111001110101;
        13: y = 16'b0010000011000010;
        14: y = 16'b0010001100000001;
        15: y = 16'b0010010100110000;
        16: y = 16'b0010011101001111;
        17: y = 16'b0010100101011100;
        18: y = 16'b0010101101011000;
        19: y = 16'b0010110101000001;
        20: y = 16'b0010111100010101;
        21: y = 16'b0011000011010110;
        22: y = 16'b0011001010000000;
        23: y = 16'b0011010000010101;
        24: y = 16'b0011010110010011;
        25: y = 16'b0011011011111010;
        26: y = 16'b0011100001001000;
        27: y = 16'b0011100101111110;
        28: y = 16'b0011101010011011;
        29: y = 16'b0011101110011110;
        30: y = 16'b0011110010000111;
        31: y = 16'b0011110101010110;
        32: y = 16'b0011111000001010;
        33: y = 16'b0011111010100010;
        34: y = 16'b0011111100100000;
        35: y = 16'b0011111110000001;
        36: y = 16'b0011111111000111;
        37: y = 16'b0011111111110001;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(pi*F*t/2), F=349.23Hz, Fs=48828Hz, 16-bit

module table_48828_F
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 34;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001011011111;
        2: y = 16'b0000010110111101;
        3: y = 16'b0000100010010111;
        4: y = 16'b0000101101101101;
        5: y = 16'b0000111000111110;
        6: y = 16'b0001000100000110;
        7: y = 16'b0001001111000111;
        8: y = 16'b0001011001111101;
        9: y = 16'b0001100100100111;
        10: y = 16'b0001101111000100;
        11: y = 16'b0001111001010011;
        12: y = 16'b0010000011010011;
        13: y = 16'b0010001101000001;
        14: y = 16'b0010010110011110;
        15: y = 16'b0010011111100111;
        16: y = 16'b0010101000011011;
        17: y = 16'b0010110000111010;
        18: y = 16'b0010111001000010;
        19: y = 16'b0011000000110010;
        20: y = 16'b0011001000001001;
        21: y = 16'b0011001111000110;
        22: y = 16'b0011010101101001;
        23: y = 16'b0011011011110000;
        24: y = 16'b0011100001011011;
        25: y = 16'b0011100110101001;
        26: y = 16'b0011101011011001;
        27: y = 16'b0011101111101010;
        28: y = 16'b0011110011011101;
        29: y = 16'b0011110110110001;
        30: y = 16'b0011111001100100;
        31: y = 16'b0011111011111000;
        32: y = 16'b0011111101101011;
        33: y = 16'b0011111110111101;
        34: y = 16'b0011111111101111;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(pi*F*t/2), F=369.99Hz, Fs=48828Hz, 16-bit

module table_48828_Fs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 32;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001100001100;
        2: y = 16'b0000011000010101;
        3: y = 16'b0000100100011100;
        4: y = 16'b0000110000011101;
        5: y = 16'b0000111100010110;
        6: y = 16'b0001001000001000;
        7: y = 16'b0001010011101110;
        8: y = 16'b0001011111001001;
        9: y = 16'b0001101010010110;
        10: y = 16'b0001110101010011;
        11: y = 16'b0001111111111111;
        12: y = 16'b0010001010011001;
        13: y = 16'b0010010100011111;
        14: y = 16'b0010011110001111;
        15: y = 16'b0010100111101001;
        16: y = 16'b0010110000101010;
        17: y = 16'b0010111001010001;
        18: y = 16'b0011000001011101;
        19: y = 16'b0011001001001110;
        20: y = 16'b0011010000100001;
        21: y = 16'b0011010111010110;
        22: y = 16'b0011011101101100;
        23: y = 16'b0011100011100010;
        24: y = 16'b0011101000110111;
        25: y = 16'b0011101101101001;
        26: y = 16'b0011110001111010;
        27: y = 16'b0011110101100111;
        28: y = 16'b0011111000110001;
        29: y = 16'b0011111011010111;
        30: y = 16'b0011111101011000;
        31: y = 16'b0011111110110101;
        32: y = 16'b0011111111101100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(pi*F*t/2), F=392.0Hz, Fs=48828Hz, 16-bit

module table_48828_G
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 31;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001100100100;
        2: y = 16'b0000011001000110;
        3: y = 16'b0000100101100100;
        4: y = 16'b0000110001111100;
        5: y = 16'b0000111110001101;
        6: y = 16'b0001001010010100;
        7: y = 16'b0001010110001111;
        8: y = 16'b0001100001111110;
        9: y = 16'b0001101101011101;
        10: y = 16'b0001111000101011;
        11: y = 16'b0010000011100111;
        12: y = 16'b0010001110001110;
        13: y = 16'b0010011000011111;
        14: y = 16'b0010100010011001;
        15: y = 16'b0010101011111010;
        16: y = 16'b0010110101000001;
        17: y = 16'b0010111101101011;
        18: y = 16'b0011000101111000;
        19: y = 16'b0011001101100111;
        20: y = 16'b0011010100110110;
        21: y = 16'b0011011011100100;
        22: y = 16'b0011100001110001;
        23: y = 16'b0011100111011010;
        24: y = 16'b0011101100100000;
        25: y = 16'b0011110001000001;
        26: y = 16'b0011110100111110;
        27: y = 16'b0011111000010100;
        28: y = 16'b0011111011000100;
        29: y = 16'b0011111101001110;
        30: y = 16'b0011111110110000;
        31: y = 16'b0011111111101011;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(pi*F*t/2), F=415.3Hz, Fs=48828Hz, 16-bit

module table_48828_Gs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 29;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001101011001;
        2: y = 16'b0000011010110000;
        3: y = 16'b0000101000000011;
        4: y = 16'b0000110101001110;
        5: y = 16'b0001000010010000;
        6: y = 16'b0001001111000111;
        7: y = 16'b0001011011101111;
        8: y = 16'b0001101000001000;
        9: y = 16'b0001110100001110;
        10: y = 16'b0001111111111111;
        11: y = 16'b0010001011011011;
        12: y = 16'b0010010110011110;
        13: y = 16'b0010100001000110;
        14: y = 16'b0010101011010010;
        15: y = 16'b0010110101000001;
        16: y = 16'b0010111110001111;
        17: y = 16'b0011000110111100;
        18: y = 16'b0011001111000110;
        19: y = 16'b0011010110101100;
        20: y = 16'b0011011101101100;
        21: y = 16'b0011100100000101;
        22: y = 16'b0011101001110111;
        23: y = 16'b0011101110111111;
        24: y = 16'b0011110011011101;
        25: y = 16'b0011110111010001;
        26: y = 16'b0011111010011001;
        27: y = 16'b0011111100110101;
        28: y = 16'b0011111110100101;
        29: y = 16'b0011111111101001;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(pi*F*t/2), F=440.0Hz, Fs=48828Hz, 16-bit

module table_48828_A
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 27;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001110010111;
        2: y = 16'b0000011100101010;
        3: y = 16'b0000101010111000;
        4: y = 16'b0000111000111110;
        5: y = 16'b0001000110110111;
        6: y = 16'b0001010100100011;
        7: y = 16'b0001100001111110;
        8: y = 16'b0001101111000100;
        9: y = 16'b0001111011110101;
        10: y = 16'b0010001000001100;
        11: y = 16'b0010010100001000;
        12: y = 16'b0010011111100111;
        13: y = 16'b0010101010100101;
        14: y = 16'b0010110101000001;
        15: y = 16'b0010111110111000;
        16: y = 16'b0011001000001001;
        17: y = 16'b0011010000110001;
        18: y = 16'b0011011000110000;
        19: y = 16'b0011100000000011;
        20: y = 16'b0011100110101001;
        21: y = 16'b0011101100100000;
        22: y = 16'b0011110001101000;
        23: y = 16'b0011110101111111;
        24: y = 16'b0011111001100100;
        25: y = 16'b0011111100011000;
        26: y = 16'b0011111110011000;
        27: y = 16'b0011111111100101;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(pi*F*t/2), F=466.16Hz, Fs=48828Hz, 16-bit

module table_48828_As
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 26;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001110111001;
        2: y = 16'b0000011101101110;
        3: y = 16'b0000101100011101;
        4: y = 16'b0000111011000010;
        5: y = 16'b0001001001011011;
        6: y = 16'b0001010111100011;
        7: y = 16'b0001100101011001;
        8: y = 16'b0001110010111001;
        9: y = 16'b0001111111111111;
        10: y = 16'b0010001100101011;
        11: y = 16'b0010011000110111;
        12: y = 16'b0010100100100011;
        13: y = 16'b0010101111101011;
        14: y = 16'b0010111010001101;
        15: y = 16'b0011000100000110;
        16: y = 16'b0011001101010101;
        17: y = 16'b0011010101111000;
        18: y = 16'b0011011101101100;
        19: y = 16'b0011100100110000;
        20: y = 16'b0011101011000011;
        21: y = 16'b0011110000100011;
        22: y = 16'b0011110101001111;
        23: y = 16'b0011111001000101;
        24: y = 16'b0011111100000110;
        25: y = 16'b0011111110010000;
        26: y = 16'b0011111111100011;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(pi*F*t/2), F=493.88Hz, Fs=48828Hz, 16-bit

module table_48828_B
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 24;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000010000000101;
        2: y = 16'b0000100000000101;
        3: y = 16'b0000101111111110;
        4: y = 16'b0000111111101010;
        5: y = 16'b0001001111000111;
        6: y = 16'b0001011110001111;
        7: y = 16'b0001101101000000;
        8: y = 16'b0001111011010101;
        9: y = 16'b0010001001001010;
        10: y = 16'b0010010110011110;
        11: y = 16'b0010100011001011;
        12: y = 16'b0010101111001111;
        13: y = 16'b0010111010100111;
        14: y = 16'b0011000101001111;
        15: y = 16'b0011001111000110;
        16: y = 16'b0011011000001001;
        17: y = 16'b0011100000010101;
        18: y = 16'b0011100111101000;
        19: y = 16'b0011101110000001;
        20: y = 16'b0011110011011101;
        21: y = 16'b0011110111111100;
        22: y = 16'b0011111011011101;
        23: y = 16'b0011111101111110;
        24: y = 16'b0011111111011111;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(pi*F*t/2), F=261.63Hz, Fs=64453Hz, 16-bit

module table_64453_C
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 61;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000000110011111;
        2: y = 16'b0000001100111110;
        3: y = 16'b0000010011011100;
        4: y = 16'b0000011001111001;
        5: y = 16'b0000100000010110;
        6: y = 16'b0000100110110001;
        7: y = 16'b0000101101001010;
        8: y = 16'b0000110011100010;
        9: y = 16'b0000111001110111;
        10: y = 16'b0001000000001010;
        11: y = 16'b0001000110011011;
        12: y = 16'b0001001100101000;
        13: y = 16'b0001010010110011;
        14: y = 16'b0001011000111010;
        15: y = 16'b0001011110111101;
        16: y = 16'b0001100100111101;
        17: y = 16'b0001101010111000;
        18: y = 16'b0001110000101111;
        19: y = 16'b0001110110100001;
        20: y = 16'b0001111100001111;
        21: y = 16'b0010000001110111;
        22: y = 16'b0010000111011010;
        23: y = 16'b0010001100110111;
        24: y = 16'b0010010010001111;
        25: y = 16'b0010010111100001;
        26: y = 16'b0010011100101100;
        27: y = 16'b0010100001110001;
        28: y = 16'b0010100110101111;
        29: y = 16'b0010101011100111;
        30: y = 16'b0010110000010111;
        31: y = 16'b0010110101000001;
        32: y = 16'b0010111001100010;
        33: y = 16'b0010111101111100;
        34: y = 16'b0011000010001111;
        35: y = 16'b0011000110011001;
        36: y = 16'b0011001010011011;
        37: y = 16'b0011001110010101;
        38: y = 16'b0011010010000111;
        39: y = 16'b0011010101101111;
        40: y = 16'b0011011001001111;
        41: y = 16'b0011011100100110;
        42: y = 16'b0011011111110100;
        43: y = 16'b0011100010111001;
        44: y = 16'b0011100101110101;
        45: y = 16'b0011101000100111;
        46: y = 16'b0011101011001111;
        47: y = 16'b0011101101101110;
        48: y = 16'b0011110000000011;
        49: y = 16'b0011110010001110;
        50: y = 16'b0011110100010000;
        51: y = 16'b0011110110000111;
        52: y = 16'b0011110111110100;
        53: y = 16'b0011111001010111;
        54: y = 16'b0011111010110000;
        55: y = 16'b0011111011111110;
        56: y = 16'b0011111101000010;
        57: y = 16'b0011111101111100;
        58: y = 16'b0011111110101011;
        59: y = 16'b0011111111010000;
        60: y = 16'b0011111111101010;
        61: y = 16'b0011111111111010;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(pi*F*t/2), F=277.18Hz, Fs=64453Hz, 16-bit

module table_64453_Cs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 58;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000000110110100;
        2: y = 16'b0000001101101000;
        3: y = 16'b0000010100011011;
        4: y = 16'b0000011011001101;
        5: y = 16'b0000100001111110;
        6: y = 16'b0000101000101110;
        7: y = 16'b0000101111011100;
        8: y = 16'b0000110110000111;
        9: y = 16'b0000111100110000;
        10: y = 16'b0001000011010110;
        11: y = 16'b0001001001111010;
        12: y = 16'b0001010000011010;
        13: y = 16'b0001010110110110;
        14: y = 16'b0001011101001110;
        15: y = 16'b0001100011100010;
        16: y = 16'b0001101001110010;
        17: y = 16'b0001101111111100;
        18: y = 16'b0001110110000010;
        19: y = 16'b0001111100000010;
        20: y = 16'b0010000001111101;
        21: y = 16'b0010000111110010;
        22: y = 16'b0010001101100001;
        23: y = 16'b0010010011001001;
        24: y = 16'b0010011000101010;
        25: y = 16'b0010011110000101;
        26: y = 16'b0010100011011000;
        27: y = 16'b0010101000100100;
        28: y = 16'b0010101101101001;
        29: y = 16'b0010110010100101;
        30: y = 16'b0010110111011010;
        31: y = 16'b0010111100000110;
        32: y = 16'b0011000000101001;
        33: y = 16'b0011000101000100;
        34: y = 16'b0011001001010110;
        35: y = 16'b0011001101011111;
        36: y = 16'b0011010001011110;
        37: y = 16'b0011010101010100;
        38: y = 16'b0011011001000000;
        39: y = 16'b0011011100100011;
        40: y = 16'b0011011111111011;
        41: y = 16'b0011100011001001;
        42: y = 16'b0011100110001101;
        43: y = 16'b0011101001000111;
        44: y = 16'b0011101011110110;
        45: y = 16'b0011101110011010;
        46: y = 16'b0011110000110011;
        47: y = 16'b0011110011000010;
        48: y = 16'b0011110101000101;
        49: y = 16'b0011110110111110;
        50: y = 16'b0011111000101011;
        51: y = 16'b0011111010001101;
        52: y = 16'b0011111011100011;
        53: y = 16'b0011111100101110;
        54: y = 16'b0011111101101110;
        55: y = 16'b0011111110100010;
        56: y = 16'b0011111111001011;
        57: y = 16'b0011111111101000;
        58: y = 16'b0011111111111001;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(pi*F*t/2), F=293.66Hz, Fs=64453Hz, 16-bit

module table_64453_D
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 54;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000000111010100;
        2: y = 16'b0000001110100111;
        3: y = 16'b0000010101111010;
        4: y = 16'b0000011101001100;
        5: y = 16'b0000100100011100;
        6: y = 16'b0000101011101010;
        7: y = 16'b0000110010110110;
        8: y = 16'b0000111001111111;
        9: y = 16'b0001000001000101;
        10: y = 16'b0001001000001000;
        11: y = 16'b0001001111000111;
        12: y = 16'b0001010110000001;
        13: y = 16'b0001011100111000;
        14: y = 16'b0001100011101001;
        15: y = 16'b0001101010010110;
        16: y = 16'b0001110000111101;
        17: y = 16'b0001110111011101;
        18: y = 16'b0001111101111000;
        19: y = 16'b0010000100001100;
        20: y = 16'b0010001010011001;
        21: y = 16'b0010010000011111;
        22: y = 16'b0010010110011110;
        23: y = 16'b0010011100010100;
        24: y = 16'b0010100010000011;
        25: y = 16'b0010100111101001;
        26: y = 16'b0010101101000110;
        27: y = 16'b0010110010011010;
        28: y = 16'b0010110111100101;
        29: y = 16'b0010111100100110;
        30: y = 16'b0011000001011101;
        31: y = 16'b0011000110001011;
        32: y = 16'b0011001010101110;
        33: y = 16'b0011001111000110;
        34: y = 16'b0011010011010100;
        35: y = 16'b0011010111010110;
        36: y = 16'b0011011011001110;
        37: y = 16'b0011011110111001;
        38: y = 16'b0011100010011010;
        39: y = 16'b0011100101101110;
        40: y = 16'b0011101000110111;
        41: y = 16'b0011101011110011;
        42: y = 16'b0011101110100011;
        43: y = 16'b0011110001000110;
        44: y = 16'b0011110011011101;
        45: y = 16'b0011110101100111;
        46: y = 16'b0011110111100101;
        47: y = 16'b0011111001010101;
        48: y = 16'b0011111010111001;
        49: y = 16'b0011111100001111;
        50: y = 16'b0011111101011000;
        51: y = 16'b0011111110010100;
        52: y = 16'b0011111111000011;
        53: y = 16'b0011111111100100;
        54: y = 16'b0011111111111000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(pi*F*t/2), F=311.13Hz, Fs=64453Hz, 16-bit

module table_64453_Ds
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 51;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000000111101111;
        2: y = 16'b0000001111011101;
        3: y = 16'b0000010111001011;
        4: y = 16'b0000011110110111;
        5: y = 16'b0000100110100001;
        6: y = 16'b0000101110001001;
        7: y = 16'b0000110101101110;
        8: y = 16'b0000111101010001;
        9: y = 16'b0001000100101111;
        10: y = 16'b0001001100001010;
        11: y = 16'b0001010011100000;
        12: y = 16'b0001011010110001;
        13: y = 16'b0001100001111110;
        14: y = 16'b0001101001000100;
        15: y = 16'b0001110000000100;
        16: y = 16'b0001110110111110;
        17: y = 16'b0001111101110000;
        18: y = 16'b0010000100011100;
        19: y = 16'b0010001010111111;
        20: y = 16'b0010010001011011;
        21: y = 16'b0010010111101110;
        22: y = 16'b0010011101111000;
        23: y = 16'b0010100011111001;
        24: y = 16'b0010101001110000;
        25: y = 16'b0010101111011101;
        26: y = 16'b0010110101000001;
        27: y = 16'b0010111010011001;
        28: y = 16'b0010111111100111;
        29: y = 16'b0011000100101001;
        30: y = 16'b0011001001100000;
        31: y = 16'b0011001110001100;
        32: y = 16'b0011010010101011;
        33: y = 16'b0011010110111110;
        34: y = 16'b0011011011000100;
        35: y = 16'b0011011110111110;
        36: y = 16'b0011100010101010;
        37: y = 16'b0011100110001010;
        38: y = 16'b0011101001011100;
        39: y = 16'b0011101100100000;
        40: y = 16'b0011101111010110;
        41: y = 16'b0011110001111111;
        42: y = 16'b0011110100011001;
        43: y = 16'b0011110110100101;
        44: y = 16'b0011111000100011;
        45: y = 16'b0011111010010010;
        46: y = 16'b0011111011110011;
        47: y = 16'b0011111101000100;
        48: y = 16'b0011111110001000;
        49: y = 16'b0011111110111100;
        50: y = 16'b0011111111100001;
        51: y = 16'b0011111111111000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(pi*F*t/2), F=329.63Hz, Fs=64453Hz, 16-bit

module table_64453_E
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 48;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001000001101;
        2: y = 16'b0000010000011010;
        3: y = 16'b0000011000100101;
        4: y = 16'b0000100000101111;
        5: y = 16'b0000101000110111;
        6: y = 16'b0000110000111100;
        7: y = 16'b0000111000111110;
        8: y = 16'b0001000000111100;
        9: y = 16'b0001001000110101;
        10: y = 16'b0001010000101010;
        11: y = 16'b0001011000011010;
        12: y = 16'b0001100000000100;
        13: y = 16'b0001100111101000;
        14: y = 16'b0001101111000100;
        15: y = 16'b0001110110011010;
        16: y = 16'b0001111101100111;
        17: y = 16'b0010000100101101;
        18: y = 16'b0010001011101001;
        19: y = 16'b0010010010011101;
        20: y = 16'b0010011001000111;
        21: y = 16'b0010011111100111;
        22: y = 16'b0010100101111100;
        23: y = 16'b0010101100000110;
        24: y = 16'b0010110010000101;
        25: y = 16'b0010110111111001;
        26: y = 16'b0010111101100000;
        27: y = 16'b0011000010111011;
        28: y = 16'b0011001000001001;
        29: y = 16'b0011001101001010;
        30: y = 16'b0011010001111101;
        31: y = 16'b0011010110100010;
        32: y = 16'b0011011010111010;
        33: y = 16'b0011011111000011;
        34: y = 16'b0011100010111101;
        35: y = 16'b0011100110101001;
        36: y = 16'b0011101010000101;
        37: y = 16'b0011101101010010;
        38: y = 16'b0011110000001111;
        39: y = 16'b0011110010111100;
        40: y = 16'b0011110101011010;
        41: y = 16'b0011110111100111;
        42: y = 16'b0011111001100100;
        43: y = 16'b0011111011010001;
        44: y = 16'b0011111100101101;
        45: y = 16'b0011111101111000;
        46: y = 16'b0011111110110011;
        47: y = 16'b0011111111011101;
        48: y = 16'b0011111111110111;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(pi*F*t/2), F=349.23Hz, Fs=64453Hz, 16-bit

module table_64453_F
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 46;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001000100011;
        2: y = 16'b0000010001000110;
        3: y = 16'b0000011001101000;
        4: y = 16'b0000100010001000;
        5: y = 16'b0000101010100101;
        6: y = 16'b0000110010111111;
        7: y = 16'b0000111011010110;
        8: y = 16'b0001000011101000;
        9: y = 16'b0001001011110110;
        10: y = 16'b0001010011111110;
        11: y = 16'b0001011100000000;
        12: y = 16'b0001100011111100;
        13: y = 16'b0001101011110000;
        14: y = 16'b0001110011011101;
        15: y = 16'b0001111011000001;
        16: y = 16'b0010000010011101;
        17: y = 16'b0010001001101111;
        18: y = 16'b0010010000111000;
        19: y = 16'b0010010111110110;
        20: y = 16'b0010011110101001;
        21: y = 16'b0010100101010001;
        22: y = 16'b0010101011101101;
        23: y = 16'b0010110001111101;
        24: y = 16'b0010111000000000;
        25: y = 16'b0010111101110110;
        26: y = 16'b0011000011011111;
        27: y = 16'b0011001000111001;
        28: y = 16'b0011001110000101;
        29: y = 16'b0011010011000011;
        30: y = 16'b0011010111110001;
        31: y = 16'b0011011100010000;
        32: y = 16'b0011100000011111;
        33: y = 16'b0011100100011110;
        34: y = 16'b0011101000001101;
        35: y = 16'b0011101011101011;
        36: y = 16'b0011101110111000;
        37: y = 16'b0011110001110101;
        38: y = 16'b0011110100011111;
        39: y = 16'b0011110110111001;
        40: y = 16'b0011111001000001;
        41: y = 16'b0011111010110111;
        42: y = 16'b0011111100011011;
        43: y = 16'b0011111101101101;
        44: y = 16'b0011111110101101;
        45: y = 16'b0011111111011010;
        46: y = 16'b0011111111110110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(pi*F*t/2), F=369.99Hz, Fs=64453Hz, 16-bit

module table_64453_Fs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 43;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001001001001;
        2: y = 16'b0000010010010001;
        3: y = 16'b0000011011010111;
        4: y = 16'b0000100100011100;
        5: y = 16'b0000101101011101;
        6: y = 16'b0000110110011010;
        7: y = 16'b0000111111010100;
        8: y = 16'b0001001000001000;
        9: y = 16'b0001010000110110;
        10: y = 16'b0001011001011101;
        11: y = 16'b0001100001111110;
        12: y = 16'b0001101010010110;
        13: y = 16'b0001110010100101;
        14: y = 16'b0001111010101100;
        15: y = 16'b0010000010101000;
        16: y = 16'b0010001010011001;
        17: y = 16'b0010010010000000;
        18: y = 16'b0010011001011010;
        19: y = 16'b0010100000101000;
        20: y = 16'b0010100111101001;
        21: y = 16'b0010101110011100;
        22: y = 16'b0010110101000001;
        23: y = 16'b0010111011010111;
        24: y = 16'b0011000001011101;
        25: y = 16'b0011000111010100;
        26: y = 16'b0011001100111011;
        27: y = 16'b0011010010010001;
        28: y = 16'b0011010111010110;
        29: y = 16'b0011011100001010;
        30: y = 16'b0011100000101011;
        31: y = 16'b0011100100111010;
        32: y = 16'b0011101000110111;
        33: y = 16'b0011101100100000;
        34: y = 16'b0011101111110110;
        35: y = 16'b0011110010111001;
        36: y = 16'b0011110101100111;
        37: y = 16'b0011111000000010;
        38: y = 16'b0011111010001001;
        39: y = 16'b0011111011111011;
        40: y = 16'b0011111101011000;
        41: y = 16'b0011111110100001;
        42: y = 16'b0011111111010101;
        43: y = 16'b0011111111110101;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(pi*F*t/2), F=392.0Hz, Fs=64453Hz, 16-bit

module table_64453_G
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 41;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001001100101;
        2: y = 16'b0000010011001000;
        3: y = 16'b0000011100101010;
        4: y = 16'b0000100110001010;
        5: y = 16'b0000101111100110;
        6: y = 16'b0000111000111110;
        7: y = 16'b0001000010010000;
        8: y = 16'b0001001011011101;
        9: y = 16'b0001010100100011;
        10: y = 16'b0001011101100001;
        11: y = 16'b0001100110010111;
        12: y = 16'b0001101111000100;
        13: y = 16'b0001110111100111;
        14: y = 16'b0001111111111111;
        15: y = 16'b0010001000001100;
        16: y = 16'b0010010000001101;
        17: y = 16'b0010011000000001;
        18: y = 16'b0010011111100111;
        19: y = 16'b0010100110111110;
        20: y = 16'b0010101110000111;
        21: y = 16'b0010110101000001;
        22: y = 16'b0010111011101010;
        23: y = 16'b0011000010000010;
        24: y = 16'b0011001000001001;
        25: y = 16'b0011001101111110;
        26: y = 16'b0011010011100000;
        27: y = 16'b0011011000110000;
        28: y = 16'b0011011101101100;
        29: y = 16'b0011100010010100;
        30: y = 16'b0011100110101001;
        31: y = 16'b0011101010101000;
        32: y = 16'b0011101110010011;
        33: y = 16'b0011110001101000;
        34: y = 16'b0011110100100111;
        35: y = 16'b0011110111010001;
        36: y = 16'b0011111001100100;
        37: y = 16'b0011111011100001;
        38: y = 16'b0011111101001000;
        39: y = 16'b0011111110011000;
        40: y = 16'b0011111111010001;
        41: y = 16'b0011111111110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(pi*F*t/2), F=415.3Hz, Fs=64453Hz, 16-bit

module table_64453_Gs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 38;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001010010100;
        2: y = 16'b0000010100100110;
        3: y = 16'b0000011110110111;
        4: y = 16'b0000101001000100;
        5: y = 16'b0000110011001101;
        6: y = 16'b0000111101010001;
        7: y = 16'b0001000111001110;
        8: y = 16'b0001010001000100;
        9: y = 16'b0001011010110001;
        10: y = 16'b0001100100010110;
        11: y = 16'b0001101101101111;
        12: y = 16'b0001110110111110;
        13: y = 16'b0010000000000000;
        14: y = 16'b0010001000110100;
        15: y = 16'b0010010001011011;
        16: y = 16'b0010011001110010;
        17: y = 16'b0010100001111001;
        18: y = 16'b0010101001110000;
        19: y = 16'b0010110001010101;
        20: y = 16'b0010111000100111;
        21: y = 16'b0010111111100111;
        22: y = 16'b0011000110010010;
        23: y = 16'b0011001100101001;
        24: y = 16'b0011010010101011;
        25: y = 16'b0011011000010111;
        26: y = 16'b0011011101101100;
        27: y = 16'b0011100010101010;
        28: y = 16'b0011100111010001;
        29: y = 16'b0011101011100000;
        30: y = 16'b0011101111010110;
        31: y = 16'b0011110010110100;
        32: y = 16'b0011110101111000;
        33: y = 16'b0011111000100011;
        34: y = 16'b0011111010110100;
        35: y = 16'b0011111100101011;
        36: y = 16'b0011111110001000;
        37: y = 16'b0011111111001010;
        38: y = 16'b0011111111110010;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(pi*F*t/2), F=440.0Hz, Fs=64453Hz, 16-bit

module table_64453_A
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 36;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001010110111;
        2: y = 16'b0000010101101101;
        3: y = 16'b0000100000100001;
        4: y = 16'b0000101011010001;
        5: y = 16'b0000110101111100;
        6: y = 16'b0001000000100000;
        7: y = 16'b0001001010111101;
        8: y = 16'b0001010101010010;
        9: y = 16'b0001011111011101;
        10: y = 16'b0001101001011100;
        11: y = 16'b0001110011010000;
        12: y = 16'b0001111100110110;
        13: y = 16'b0010000110001110;
        14: y = 16'b0010001111010110;
        15: y = 16'b0010011000001110;
        16: y = 16'b0010100000110100;
        17: y = 16'b0010101001001000;
        18: y = 16'b0010110001001000;
        19: y = 16'b0010111000110100;
        20: y = 16'b0011000000001010;
        21: y = 16'b0011000111001011;
        22: y = 16'b0011001101110100;
        23: y = 16'b0011010100000101;
        24: y = 16'b0011011001111111;
        25: y = 16'b0011011111011111;
        26: y = 16'b0011100100100101;
        27: y = 16'b0011101001010001;
        28: y = 16'b0011101101100010;
        29: y = 16'b0011110001010111;
        30: y = 16'b0011110100110001;
        31: y = 16'b0011110111101110;
        32: y = 16'b0011111010001111;
        33: y = 16'b0011111100010011;
        34: y = 16'b0011111101111010;
        35: y = 16'b0011111111000100;
        36: y = 16'b0011111111110000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(pi*F*t/2), F=466.16Hz, Fs=64453Hz, 16-bit

module table_64453_As
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 34;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001011011111;
        2: y = 16'b0000010110111101;
        3: y = 16'b0000100010010111;
        4: y = 16'b0000101101101101;
        5: y = 16'b0000111000111110;
        6: y = 16'b0001000100000110;
        7: y = 16'b0001001111000111;
        8: y = 16'b0001011001111101;
        9: y = 16'b0001100100100111;
        10: y = 16'b0001101111000100;
        11: y = 16'b0001111001010011;
        12: y = 16'b0010000011010011;
        13: y = 16'b0010001101000001;
        14: y = 16'b0010010110011110;
        15: y = 16'b0010011111100111;
        16: y = 16'b0010101000011011;
        17: y = 16'b0010110000111010;
        18: y = 16'b0010111001000010;
        19: y = 16'b0011000000110010;
        20: y = 16'b0011001000001001;
        21: y = 16'b0011001111000110;
        22: y = 16'b0011010101101001;
        23: y = 16'b0011011011110000;
        24: y = 16'b0011100001011011;
        25: y = 16'b0011100110101001;
        26: y = 16'b0011101011011001;
        27: y = 16'b0011101111101010;
        28: y = 16'b0011110011011101;
        29: y = 16'b0011110110110001;
        30: y = 16'b0011111001100100;
        31: y = 16'b0011111011111000;
        32: y = 16'b0011111101101011;
        33: y = 16'b0011111110111101;
        34: y = 16'b0011111111101111;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(pi*F*t/2), F=493.88Hz, Fs=64453Hz, 16-bit

module table_64453_B
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 32;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001100001100;
        2: y = 16'b0000011000010101;
        3: y = 16'b0000100100011100;
        4: y = 16'b0000110000011101;
        5: y = 16'b0000111100010110;
        6: y = 16'b0001001000001000;
        7: y = 16'b0001010011101110;
        8: y = 16'b0001011111001001;
        9: y = 16'b0001101010010110;
        10: y = 16'b0001110101010011;
        11: y = 16'b0001111111111111;
        12: y = 16'b0010001010011001;
        13: y = 16'b0010010100011111;
        14: y = 16'b0010011110001111;
        15: y = 16'b0010100111101001;
        16: y = 16'b0010110000101010;
        17: y = 16'b0010111001010001;
        18: y = 16'b0011000001011101;
        19: y = 16'b0011001001001110;
        20: y = 16'b0011010000100001;
        21: y = 16'b0011010111010110;
        22: y = 16'b0011011101101100;
        23: y = 16'b0011100011100010;
        24: y = 16'b0011101000110111;
        25: y = 16'b0011101101101001;
        26: y = 16'b0011110001111010;
        27: y = 16'b0011110101100111;
        28: y = 16'b0011111000110001;
        29: y = 16'b0011111011010111;
        30: y = 16'b0011111101011000;
        31: y = 16'b0011111110110101;
        32: y = 16'b0011111111101100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(pi*F*t/2), F=261.63Hz, Fs=52734Hz, 16-bit

module table_52734_C
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 50;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000000111111001;
        2: y = 16'b0000001111110001;
        3: y = 16'b0000010111101000;
        4: y = 16'b0000011111011101;
        5: y = 16'b0000100111010001;
        6: y = 16'b0000101111000010;
        7: y = 16'b0000110110110001;
        8: y = 16'b0000111110011100;
        9: y = 16'b0001000110000011;
        10: y = 16'b0001001101100111;
        11: y = 16'b0001010101000101;
        12: y = 16'b0001011100011110;
        13: y = 16'b0001100011110010;
        14: y = 16'b0001101010111111;
        15: y = 16'b0001110010000111;
        16: y = 16'b0001111001000111;
        17: y = 16'b0010000000000000;
        18: y = 16'b0010000110110001;
        19: y = 16'b0010001101011001;
        20: y = 16'b0010010011111010;
        21: y = 16'b0010011010010001;
        22: y = 16'b0010100000011111;
        23: y = 16'b0010100110100011;
        24: y = 16'b0010101100011101;
        25: y = 16'b0010110010001101;
        26: y = 16'b0010110111110010;
        27: y = 16'b0010111101001011;
        28: y = 16'b0011000010011001;
        29: y = 16'b0011000111011100;
        30: y = 16'b0011001100010010;
        31: y = 16'b0011010000111100;
        32: y = 16'b0011010101011001;
        33: y = 16'b0011011001101001;
        34: y = 16'b0011011101101100;
        35: y = 16'b0011100001100010;
        36: y = 16'b0011100101001001;
        37: y = 16'b0011101000100011;
        38: y = 16'b0011101011101111;
        39: y = 16'b0011101110101101;
        40: y = 16'b0011110001011100;
        41: y = 16'b0011110011111100;
        42: y = 16'b0011110110001110;
        43: y = 16'b0011111000010000;
        44: y = 16'b0011111010000100;
        45: y = 16'b0011111011101000;
        46: y = 16'b0011111100111101;
        47: y = 16'b0011111110000011;
        48: y = 16'b0011111110111001;
        49: y = 16'b0011111111100000;
        50: y = 16'b0011111111110111;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(pi*F*t/2), F=277.18Hz, Fs=52734Hz, 16-bit

module table_52734_Cs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 47;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001000011000;
        2: y = 16'b0000010000101111;
        3: y = 16'b0000011001000110;
        4: y = 16'b0000100001011010;
        5: y = 16'b0000101001101101;
        6: y = 16'b0000110001111100;
        7: y = 16'b0000111010001000;
        8: y = 16'b0001000010010000;
        9: y = 16'b0001001010010100;
        10: y = 16'b0001010010010010;
        11: y = 16'b0001011010001011;
        12: y = 16'b0001100001111110;
        13: y = 16'b0001101001101001;
        14: y = 16'b0001110001001110;
        15: y = 16'b0001111000101011;
        16: y = 16'b0001111111111111;
        17: y = 16'b0010000111001011;
        18: y = 16'b0010001110001110;
        19: y = 16'b0010010101000111;
        20: y = 16'b0010011011110101;
        21: y = 16'b0010100010011001;
        22: y = 16'b0010101000110010;
        23: y = 16'b0010101110111111;
        24: y = 16'b0010110101000001;
        25: y = 16'b0010111010110101;
        26: y = 16'b0011000000011101;
        27: y = 16'b0011000101111000;
        28: y = 16'b0011001011000110;
        29: y = 16'b0011010000000101;
        30: y = 16'b0011010100110110;
        31: y = 16'b0011011001011000;
        32: y = 16'b0011011101101100;
        33: y = 16'b0011100001110001;
        34: y = 16'b0011100101100101;
        35: y = 16'b0011101001001011;
        36: y = 16'b0011101100100000;
        37: y = 16'b0011101111100101;
        38: y = 16'b0011110010011010;
        39: y = 16'b0011110100111110;
        40: y = 16'b0011110111010001;
        41: y = 16'b0011111001010011;
        42: y = 16'b0011111011000100;
        43: y = 16'b0011111100100100;
        44: y = 16'b0011111101110011;
        45: y = 16'b0011111110110000;
        46: y = 16'b0011111111011100;
        47: y = 16'b0011111111110110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(pi*F*t/2), F=293.66Hz, Fs=52734Hz, 16-bit

module table_52734_D
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 44;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001000111100;
        2: y = 16'b0000010001110111;
        3: y = 16'b0000011010110000;
        4: y = 16'b0000100011101000;
        5: y = 16'b0000101100011101;
        6: y = 16'b0000110101001110;
        7: y = 16'b0000111101111011;
        8: y = 16'b0001000110100100;
        9: y = 16'b0001001111000111;
        10: y = 16'b0001010111100011;
        11: y = 16'b0001011111111001;
        12: y = 16'b0001101000001000;
        13: y = 16'b0001110000001110;
        14: y = 16'b0001111000001011;
        15: y = 16'b0001111111111111;
        16: y = 16'b0010000111101010;
        17: y = 16'b0010001111001001;
        18: y = 16'b0010010110011110;
        19: y = 16'b0010011101100110;
        20: y = 16'b0010100100100011;
        21: y = 16'b0010101011010010;
        22: y = 16'b0010110001110101;
        23: y = 16'b0010111000001001;
        24: y = 16'b0010111110001111;
        25: y = 16'b0011000100000110;
        26: y = 16'b0011001001101110;
        27: y = 16'b0011001111000110;
        28: y = 16'b0011010100001110;
        29: y = 16'b0011011001000110;
        30: y = 16'b0011011101101100;
        31: y = 16'b0011100010000001;
        32: y = 16'b0011100110000101;
        33: y = 16'b0011101001110111;
        34: y = 16'b0011101101010110;
        35: y = 16'b0011110000100011;
        36: y = 16'b0011110011011101;
        37: y = 16'b0011110110000100;
        38: y = 16'b0011111000011000;
        39: y = 16'b0011111010011001;
        40: y = 16'b0011111100000110;
        41: y = 16'b0011111101100000;
        42: y = 16'b0011111110100101;
        43: y = 16'b0011111111010111;
        44: y = 16'b0011111111110101;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(pi*F*t/2), F=311.13Hz, Fs=52734Hz, 16-bit

module table_52734_Ds
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 42;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001001010110;
        2: y = 16'b0000010010101100;
        3: y = 16'b0000011100000000;
        4: y = 16'b0000100101010001;
        5: y = 16'b0000101110100000;
        6: y = 16'b0000110111101010;
        7: y = 16'b0001000000110000;
        8: y = 16'b0001001001110000;
        9: y = 16'b0001010010101010;
        10: y = 16'b0001011011011101;
        11: y = 16'b0001100100000111;
        12: y = 16'b0001101100101010;
        13: y = 16'b0001110101000011;
        14: y = 16'b0001111101010010;
        15: y = 16'b0010000101010111;
        16: y = 16'b0010001101010000;
        17: y = 16'b0010010100111101;
        18: y = 16'b0010011100011101;
        19: y = 16'b0010100011110000;
        20: y = 16'b0010101010110101;
        21: y = 16'b0010110001101011;
        22: y = 16'b0010111000010010;
        23: y = 16'b0010111110101010;
        24: y = 16'b0011000100110001;
        25: y = 16'b0011001010100111;
        26: y = 16'b0011010000001100;
        27: y = 16'b0011010101011111;
        28: y = 16'b0011011010100000;
        29: y = 16'b0011011111001111;
        30: y = 16'b0011100011101010;
        31: y = 16'b0011100111110010;
        32: y = 16'b0011101011100110;
        33: y = 16'b0011101111000110;
        34: y = 16'b0011110010010010;
        35: y = 16'b0011110101001000;
        36: y = 16'b0011110111101010;
        37: y = 16'b0011111001110111;
        38: y = 16'b0011111011101110;
        39: y = 16'b0011111101010000;
        40: y = 16'b0011111110011101;
        41: y = 16'b0011111111010011;
        42: y = 16'b0011111111110100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(pi*F*t/2), F=329.63Hz, Fs=52734Hz, 16-bit

module table_52734_E
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 39;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001010000011;
        2: y = 16'b0000010100000101;
        3: y = 16'b0000011110000110;
        4: y = 16'b0000101000000011;
        5: y = 16'b0000110001111100;
        6: y = 16'b0000111011110001;
        7: y = 16'b0001000101011111;
        8: y = 16'b0001001111000111;
        9: y = 16'b0001011000100110;
        10: y = 16'b0001100001111110;
        11: y = 16'b0001101011001011;
        12: y = 16'b0001110100001110;
        13: y = 16'b0001111101000101;
        14: y = 16'b0010000101110000;
        15: y = 16'b0010001110001110;
        16: y = 16'b0010010110011110;
        17: y = 16'b0010011110011111;
        18: y = 16'b0010100110010000;
        19: y = 16'b0010101101110001;
        20: y = 16'b0010110101000001;
        21: y = 16'b0010111011111110;
        22: y = 16'b0011000010101010;
        23: y = 16'b0011001001000010;
        24: y = 16'b0011001111000110;
        25: y = 16'b0011010100110110;
        26: y = 16'b0011011010010001;
        27: y = 16'b0011011111010110;
        28: y = 16'b0011100100000101;
        29: y = 16'b0011101000011110;
        30: y = 16'b0011101100100000;
        31: y = 16'b0011110000001010;
        32: y = 16'b0011110011011101;
        33: y = 16'b0011110110011000;
        34: y = 16'b0011111000111010;
        35: y = 16'b0011111011000100;
        36: y = 16'b0011111100110101;
        37: y = 16'b0011111110001101;
        38: y = 16'b0011111111001100;
        39: y = 16'b0011111111110010;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(pi*F*t/2), F=349.23Hz, Fs=52734Hz, 16-bit

module table_52734_F
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 37;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001010100101;
        2: y = 16'b0000010101001001;
        3: y = 16'b0000011111101010;
        4: y = 16'b0000101010001001;
        5: y = 16'b0000110100100010;
        6: y = 16'b0000111110110110;
        7: y = 16'b0001001001000011;
        8: y = 16'b0001010011001000;
        9: y = 16'b0001011101000011;
        10: y = 16'b0001100110110101;
        11: y = 16'b0001110000011011;
        12: y = 16'b0001111001110101;
        13: y = 16'b0010000011000010;
        14: y = 16'b0010001100000001;
        15: y = 16'b0010010100110000;
        16: y = 16'b0010011101001111;
        17: y = 16'b0010100101011100;
        18: y = 16'b0010101101011000;
        19: y = 16'b0010110101000001;
        20: y = 16'b0010111100010101;
        21: y = 16'b0011000011010110;
        22: y = 16'b0011001010000000;
        23: y = 16'b0011010000010101;
        24: y = 16'b0011010110010011;
        25: y = 16'b0011011011111010;
        26: y = 16'b0011100001001000;
        27: y = 16'b0011100101111110;
        28: y = 16'b0011101010011011;
        29: y = 16'b0011101110011110;
        30: y = 16'b0011110010000111;
        31: y = 16'b0011110101010110;
        32: y = 16'b0011111000001010;
        33: y = 16'b0011111010100010;
        34: y = 16'b0011111100100000;
        35: y = 16'b0011111110000001;
        36: y = 16'b0011111111000111;
        37: y = 16'b0011111111110001;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(pi*F*t/2), F=369.99Hz, Fs=52734Hz, 16-bit

module table_52734_Fs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 35;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001011001011;
        2: y = 16'b0000010110010100;
        3: y = 16'b0000100001011010;
        4: y = 16'b0000101100011101;
        5: y = 16'b0000110111011010;
        6: y = 16'b0001000010010000;
        7: y = 16'b0001001100111110;
        8: y = 16'b0001010111100011;
        9: y = 16'b0001100001111110;
        10: y = 16'b0001101100001100;
        11: y = 16'b0001110110001101;
        12: y = 16'b0001111111111111;
        13: y = 16'b0010001001100011;
        14: y = 16'b0010010010110101;
        15: y = 16'b0010011011110101;
        16: y = 16'b0010100100100011;
        17: y = 16'b0010101100111100;
        18: y = 16'b0010110101000001;
        19: y = 16'b0010111100101111;
        20: y = 16'b0011000100000110;
        21: y = 16'b0011001011000110;
        22: y = 16'b0011010001101100;
        23: y = 16'b0011010111111001;
        24: y = 16'b0011011101101100;
        25: y = 16'b0011100011000100;
        26: y = 16'b0011101000000000;
        27: y = 16'b0011101100100000;
        28: y = 16'b0011110000100011;
        29: y = 16'b0011110100001001;
        30: y = 16'b0011110111010001;
        31: y = 16'b0011111001111011;
        32: y = 16'b0011111100000110;
        33: y = 16'b0011111101110011;
        34: y = 16'b0011111111000001;
        35: y = 16'b0011111111101111;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(pi*F*t/2), F=392.0Hz, Fs=52734Hz, 16-bit

module table_52734_G
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 33;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001011110101;
        2: y = 16'b0000010111101000;
        3: y = 16'b0000100011010111;
        4: y = 16'b0000101111000010;
        5: y = 16'b0000111010100111;
        6: y = 16'b0001000110000011;
        7: y = 16'b0001010001010110;
        8: y = 16'b0001011100011110;
        9: y = 16'b0001100111011001;
        10: y = 16'b0001110010000111;
        11: y = 16'b0001111100100100;
        12: y = 16'b0010000110110001;
        13: y = 16'b0010010000101011;
        14: y = 16'b0010011010010001;
        15: y = 16'b0010100011100010;
        16: y = 16'b0010101100011101;
        17: y = 16'b0010110101000001;
        18: y = 16'b0010111101001011;
        19: y = 16'b0011000100111100;
        20: y = 16'b0011001100010010;
        21: y = 16'b0011010011001100;
        22: y = 16'b0011011001101001;
        23: y = 16'b0011011111101001;
        24: y = 16'b0011100101001001;
        25: y = 16'b0011101010001011;
        26: y = 16'b0011101110101101;
        27: y = 16'b0011110010101110;
        28: y = 16'b0011110110001110;
        29: y = 16'b0011111001001100;
        30: y = 16'b0011111011101000;
        31: y = 16'b0011111101100010;
        32: y = 16'b0011111110111001;
        33: y = 16'b0011111111101110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(pi*F*t/2), F=415.3Hz, Fs=52734Hz, 16-bit

module table_52734_Gs
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 31;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001100100100;
        2: y = 16'b0000011001000110;
        3: y = 16'b0000100101100100;
        4: y = 16'b0000110001111100;
        5: y = 16'b0000111110001101;
        6: y = 16'b0001001010010100;
        7: y = 16'b0001010110001111;
        8: y = 16'b0001100001111110;
        9: y = 16'b0001101101011101;
        10: y = 16'b0001111000101011;
        11: y = 16'b0010000011100111;
        12: y = 16'b0010001110001110;
        13: y = 16'b0010011000011111;
        14: y = 16'b0010100010011001;
        15: y = 16'b0010101011111010;
        16: y = 16'b0010110101000001;
        17: y = 16'b0010111101101011;
        18: y = 16'b0011000101111000;
        19: y = 16'b0011001101100111;
        20: y = 16'b0011010100110110;
        21: y = 16'b0011011011100100;
        22: y = 16'b0011100001110001;
        23: y = 16'b0011100111011010;
        24: y = 16'b0011101100100000;
        25: y = 16'b0011110001000001;
        26: y = 16'b0011110100111110;
        27: y = 16'b0011111000010100;
        28: y = 16'b0011111011000100;
        29: y = 16'b0011111101001110;
        30: y = 16'b0011111110110000;
        31: y = 16'b0011111111101011;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(pi*F*t/2), F=440.0Hz, Fs=52734Hz, 16-bit

module table_52734_A
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 29;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001101011001;
        2: y = 16'b0000011010110000;
        3: y = 16'b0000101000000011;
        4: y = 16'b0000110101001110;
        5: y = 16'b0001000010010000;
        6: y = 16'b0001001111000111;
        7: y = 16'b0001011011101111;
        8: y = 16'b0001101000001000;
        9: y = 16'b0001110100001110;
        10: y = 16'b0001111111111111;
        11: y = 16'b0010001011011011;
        12: y = 16'b0010010110011110;
        13: y = 16'b0010100001000110;
        14: y = 16'b0010101011010010;
        15: y = 16'b0010110101000001;
        16: y = 16'b0010111110001111;
        17: y = 16'b0011000110111100;
        18: y = 16'b0011001111000110;
        19: y = 16'b0011010110101100;
        20: y = 16'b0011011101101100;
        21: y = 16'b0011100100000101;
        22: y = 16'b0011101001110111;
        23: y = 16'b0011101110111111;
        24: y = 16'b0011110011011101;
        25: y = 16'b0011110111010001;
        26: y = 16'b0011111010011001;
        27: y = 16'b0011111100110101;
        28: y = 16'b0011111110100101;
        29: y = 16'b0011111111101001;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(pi*F*t/2), F=466.16Hz, Fs=52734Hz, 16-bit

module table_52734_As
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 28;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001101110111;
        2: y = 16'b0000011011101011;
        3: y = 16'b0000101001011010;
        4: y = 16'b0000110111000010;
        5: y = 16'b0001000100011111;
        6: y = 16'b0001010001101111;
        7: y = 16'b0001011110110000;
        8: y = 16'b0001101011011111;
        9: y = 16'b0001110111111010;
        10: y = 16'b0010000011111110;
        11: y = 16'b0010001111101010;
        12: y = 16'b0010011010111011;
        13: y = 16'b0010100101101110;
        14: y = 16'b0010110000000011;
        15: y = 16'b0010111001110110;
        16: y = 16'b0011000011000111;
        17: y = 16'b0011001011110010;
        18: y = 16'b0011010011111000;
        19: y = 16'b0011011011010110;
        20: y = 16'b0011100010001011;
        21: y = 16'b0011101000010101;
        22: y = 16'b0011101101110011;
        23: y = 16'b0011110010100101;
        24: y = 16'b0011110110101010;
        25: y = 16'b0011111010000000;
        26: y = 16'b0011111100100111;
        27: y = 16'b0011111110011111;
        28: y = 16'b0011111111100111;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(pi*F*t/2), F=493.88Hz, Fs=52734Hz, 16-bit

module table_52734_B
(
    input        [ 8:0] x,
    output       [ 8:0] x_max,
    output logic [15:0] y
);

    assign x_max = 26;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000001110111001;
        2: y = 16'b0000011101101110;
        3: y = 16'b0000101100011101;
        4: y = 16'b0000111011000010;
        5: y = 16'b0001001001011011;
        6: y = 16'b0001010111100011;
        7: y = 16'b0001100101011001;
        8: y = 16'b0001110010111001;
        9: y = 16'b0001111111111111;
        10: y = 16'b0010001100101011;
        11: y = 16'b0010011000110111;
        12: y = 16'b0010100100100011;
        13: y = 16'b0010101111101011;
        14: y = 16'b0010111010001101;
        15: y = 16'b0011000100000110;
        16: y = 16'b0011001101010101;
        17: y = 16'b0011010101111000;
        18: y = 16'b0011011101101100;
        19: y = 16'b0011100100110000;
        20: y = 16'b0011101011000011;
        21: y = 16'b0011110000100011;
        22: y = 16'b0011110101001111;
        23: y = 16'b0011111001000101;
        24: y = 16'b0011111100000110;
        25: y = 16'b0011111110010000;
        26: y = 16'b0011111111100011;
        default: y = 16'b0;
        endcase

endmodule

